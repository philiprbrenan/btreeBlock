//-----------------------------------------------------------------------------
// Generic cpu
// Philip R Brenan at appaapps dot com, Appa Apps Ltd Inc., 2025-01-07
//------------------------------------------------------------------------------
`timescale 10ps/1ps
(* keep_hierarchy = "yes" *)
module put(reset, stop, clock, Key, Data, data, found);                    // Database on a chip
  input                      reset;                                             // Restart the program run sequence when this goes high
  input                      clock;                                             // Program counter clock
  input [16-1:0]  Key;                                             // Input key
  input [16-1:0] Data;                                             // Input data
  output                      stop;                                             // Program has stopped when this goes high
  output[16-1:0] data;                                             // Output data
  output                     found;                                             // Whether the key was found on put, find delete

  integer step;
  integer steps;
  integer stopped;
  integer intermediateValue;
  reg [16-1:0] memory [351-1: 0]; /* declareVerilogMemory */
  reg [10-1: 0] opCodes[3072 : 0];

  assign stop  = stopped > 0 ? 1 : 0;
  assign found = memory[108];  // found
  assign data  = memory[107];   // data

  always @ (posedge clock) begin                                                // Execute next step in program
    if (reset) begin                                                            // Reset
      step     <= 0;
      steps    <= 0;
      stopped  <= 0;
      begin /* initilizeVerilogMemory */
        integer i;
        for (i = 0; i < 351; i = i + 1) begin
          memory[i] <= 0;
        end
      end
      memory[ 119] <=    1; /* freeChainHead */
      memory[ 121] <=    2; /* free[1] */
      memory[ 122] <=    3; /* free[2] */
      memory[ 123] <=    4; /* free[3] */
      memory[ 124] <=    5; /* free[4] */
      memory[ 125] <=    6; /* free[5] */
      memory[ 126] <=    7; /* free[6] */
      memory[ 127] <=    8; /* free[7] */
      memory[ 128] <=    9; /* free[8] */
      memory[ 129] <=   10; /* free[9] */
      memory[ 130] <=   11; /* free[10] */
      memory[ 131] <=   12; /* free[11] */
      memory[ 132] <=   13; /* free[12] */
      memory[ 133] <=   14; /* free[13] */
      memory[ 134] <=   15; /* free[14] */
      memory[ 135] <=   16; /* free[15] */
      memory[ 136] <=   17; /* free[16] */
      memory[ 137] <=   18; /* free[17] */
      memory[ 138] <=   19; /* free[18] */
      memory[ 145] <=    1; /* isLeaf[0] */

      opCodes[0] <= 0;
      opCodes[908] <= 0;
      opCodes[1303] <= 0;
      opCodes[3030] <= 0;
      opCodes[1] <= 1;
      opCodes[2] <= 2;
      opCodes[3] <= 3;
      opCodes[4] <= 4;
      opCodes[137] <= 4;
      opCodes[169] <= 4;
      opCodes[193] <= 4;
      opCodes[674] <= 4;
      opCodes[807] <= 4;
      opCodes[839] <= 4;
      opCodes[863] <= 4;
      opCodes[1076] <= 4;
      opCodes[1209] <= 4;
      opCodes[1241] <= 4;
      opCodes[1265] <= 4;
      opCodes[5] <= 5;
      opCodes[675] <= 5;
      opCodes[1077] <= 5;
      opCodes[6] <= 6;
      opCodes[264] <= 6;
      opCodes[676] <= 6;
      opCodes[1078] <= 6;
      opCodes[1305] <= 6;
      opCodes[7] <= 7;
      opCodes[265] <= 7;
      opCodes[677] <= 7;
      opCodes[1079] <= 7;
      opCodes[1306] <= 7;
      opCodes[8] <= 8;
      opCodes[266] <= 8;
      opCodes[443] <= 8;
      opCodes[678] <= 8;
      opCodes[1080] <= 8;
      opCodes[1307] <= 8;
      opCodes[9] <= 9;
      opCodes[10] <= 10;
      opCodes[680] <= 10;
      opCodes[1082] <= 10;
      opCodes[1320] <= 10;
      opCodes[11] <= 11;
      opCodes[49] <= 11;
      opCodes[88] <= 11;
      opCodes[681] <= 11;
      opCodes[719] <= 11;
      opCodes[758] <= 11;
      opCodes[1083] <= 11;
      opCodes[1121] <= 11;
      opCodes[1160] <= 11;
      opCodes[12] <= 12;
      opCodes[23] <= 12;
      opCodes[50] <= 12;
      opCodes[64] <= 12;
      opCodes[75] <= 12;
      opCodes[89] <= 12;
      opCodes[100] <= 12;
      opCodes[138] <= 12;
      opCodes[170] <= 12;
      opCodes[181] <= 12;
      opCodes[194] <= 12;
      opCodes[314] <= 12;
      opCodes[352] <= 12;
      opCodes[388] <= 12;
      opCodes[401] <= 12;
      opCodes[418] <= 12;
      opCodes[431] <= 12;
      opCodes[491] <= 12;
      opCodes[529] <= 12;
      opCodes[557] <= 12;
      opCodes[571] <= 12;
      opCodes[609] <= 12;
      opCodes[635] <= 12;
      opCodes[649] <= 12;
      opCodes[662] <= 12;
      opCodes[682] <= 12;
      opCodes[693] <= 12;
      opCodes[720] <= 12;
      opCodes[734] <= 12;
      opCodes[745] <= 12;
      opCodes[759] <= 12;
      opCodes[770] <= 12;
      opCodes[808] <= 12;
      opCodes[840] <= 12;
      opCodes[851] <= 12;
      opCodes[864] <= 12;
      opCodes[909] <= 12;
      opCodes[923] <= 12;
      opCodes[934] <= 12;
      opCodes[976] <= 12;
      opCodes[1014] <= 12;
      opCodes[1027] <= 12;
      opCodes[1042] <= 12;
      opCodes[1084] <= 12;
      opCodes[1095] <= 12;
      opCodes[1122] <= 12;
      opCodes[1136] <= 12;
      opCodes[1147] <= 12;
      opCodes[1161] <= 12;
      opCodes[1172] <= 12;
      opCodes[1210] <= 12;
      opCodes[1242] <= 12;
      opCodes[1253] <= 12;
      opCodes[1266] <= 12;
      opCodes[1323] <= 12;
      opCodes[1334] <= 12;
      opCodes[1378] <= 12;
      opCodes[1419] <= 12;
      opCodes[1460] <= 12;
      opCodes[1501] <= 12;
      opCodes[1604] <= 12;
      opCodes[1617] <= 12;
      opCodes[1658] <= 12;
      opCodes[1699] <= 12;
      opCodes[1741] <= 12;
      opCodes[1747] <= 12;
      opCodes[1764] <= 12;
      opCodes[1805] <= 12;
      opCodes[1846] <= 12;
      opCodes[1888] <= 12;
      opCodes[1894] <= 12;
      opCodes[1987] <= 12;
      opCodes[1995] <= 12;
      opCodes[2042] <= 12;
      opCodes[2083] <= 12;
      opCodes[2151] <= 12;
      opCodes[2164] <= 12;
      opCodes[2170] <= 12;
      opCodes[2204] <= 12;
      opCodes[2230] <= 12;
      opCodes[2271] <= 12;
      opCodes[2312] <= 12;
      opCodes[2375] <= 12;
      opCodes[2417] <= 12;
      opCodes[2428] <= 12;
      opCodes[2471] <= 12;
      opCodes[2512] <= 12;
      opCodes[2584] <= 12;
      opCodes[2594] <= 12;
      opCodes[2624] <= 12;
      opCodes[2665] <= 12;
      opCodes[2706] <= 12;
      opCodes[2764] <= 12;
      opCodes[2772] <= 12;
      opCodes[2776] <= 12;
      opCodes[2803] <= 12;
      opCodes[2830] <= 12;
      opCodes[2844] <= 12;
      opCodes[2855] <= 12;
      opCodes[2915] <= 12;
      opCodes[2953] <= 12;
      opCodes[2981] <= 12;
      opCodes[2994] <= 12;
      opCodes[3031] <= 12;
      opCodes[3045] <= 12;
      opCodes[3056] <= 12;
      opCodes[13] <= 13;
      opCodes[51] <= 13;
      opCodes[90] <= 13;
      opCodes[171] <= 13;
      opCodes[683] <= 13;
      opCodes[721] <= 13;
      opCodes[760] <= 13;
      opCodes[841] <= 13;
      opCodes[910] <= 13;
      opCodes[1085] <= 13;
      opCodes[1123] <= 13;
      opCodes[1162] <= 13;
      opCodes[1243] <= 13;
      opCodes[2831] <= 13;
      opCodes[3032] <= 13;
      opCodes[14] <= 14;
      opCodes[52] <= 14;
      opCodes[91] <= 14;
      opCodes[172] <= 14;
      opCodes[386] <= 14;
      opCodes[684] <= 14;
      opCodes[722] <= 14;
      opCodes[761] <= 14;
      opCodes[842] <= 14;
      opCodes[911] <= 14;
      opCodes[1012] <= 14;
      opCodes[1086] <= 14;
      opCodes[1124] <= 14;
      opCodes[1163] <= 14;
      opCodes[1244] <= 14;
      opCodes[1321] <= 14;
      opCodes[1602] <= 14;
      opCodes[2064] <= 14;
      opCodes[2105] <= 14;
      opCodes[2188] <= 14;
      opCodes[2252] <= 14;
      opCodes[2293] <= 14;
      opCodes[2334] <= 14;
      opCodes[2832] <= 14;
      opCodes[3033] <= 14;
      opCodes[15] <= 15;
      opCodes[53] <= 15;
      opCodes[92] <= 15;
      opCodes[149] <= 15;
      opCodes[173] <= 15;
      opCodes[199] <= 15;
      opCodes[223] <= 15;
      opCodes[317] <= 15;
      opCodes[334] <= 15;
      opCodes[339] <= 15;
      opCodes[345] <= 15;
      opCodes[355] <= 15;
      opCodes[372] <= 15;
      opCodes[377] <= 15;
      opCodes[383] <= 15;
      opCodes[395] <= 15;
      opCodes[421] <= 15;
      opCodes[427] <= 15;
      opCodes[434] <= 15;
      opCodes[440] <= 15;
      opCodes[494] <= 15;
      opCodes[511] <= 15;
      opCodes[516] <= 15;
      opCodes[522] <= 15;
      opCodes[532] <= 15;
      opCodes[549] <= 15;
      opCodes[558] <= 15;
      opCodes[564] <= 15;
      opCodes[574] <= 15;
      opCodes[591] <= 15;
      opCodes[596] <= 15;
      opCodes[602] <= 15;
      opCodes[612] <= 15;
      opCodes[629] <= 15;
      opCodes[636] <= 15;
      opCodes[642] <= 15;
      opCodes[652] <= 15;
      opCodes[658] <= 15;
      opCodes[665] <= 15;
      opCodes[671] <= 15;
      opCodes[685] <= 15;
      opCodes[723] <= 15;
      opCodes[762] <= 15;
      opCodes[819] <= 15;
      opCodes[843] <= 15;
      opCodes[869] <= 15;
      opCodes[893] <= 15;
      opCodes[912] <= 15;
      opCodes[979] <= 15;
      opCodes[996] <= 15;
      opCodes[1001] <= 15;
      opCodes[1007] <= 15;
      opCodes[1021] <= 15;
      opCodes[1049] <= 15;
      opCodes[1073] <= 15;
      opCodes[1087] <= 15;
      opCodes[1125] <= 15;
      opCodes[1164] <= 15;
      opCodes[1221] <= 15;
      opCodes[1245] <= 15;
      opCodes[1271] <= 15;
      opCodes[1295] <= 15;
      opCodes[1328] <= 15;
      opCodes[1381] <= 15;
      opCodes[1398] <= 15;
      opCodes[1403] <= 15;
      opCodes[1409] <= 15;
      opCodes[1422] <= 15;
      opCodes[1439] <= 15;
      opCodes[1444] <= 15;
      opCodes[1450] <= 15;
      opCodes[1463] <= 15;
      opCodes[1480] <= 15;
      opCodes[1485] <= 15;
      opCodes[1491] <= 15;
      opCodes[1504] <= 15;
      opCodes[1521] <= 15;
      opCodes[1526] <= 15;
      opCodes[1532] <= 15;
      opCodes[1620] <= 15;
      opCodes[1637] <= 15;
      opCodes[1642] <= 15;
      opCodes[1648] <= 15;
      opCodes[1661] <= 15;
      opCodes[1678] <= 15;
      opCodes[1683] <= 15;
      opCodes[1689] <= 15;
      opCodes[1702] <= 15;
      opCodes[1719] <= 15;
      opCodes[1724] <= 15;
      opCodes[1730] <= 15;
      opCodes[1735] <= 15;
      opCodes[1748] <= 15;
      opCodes[1754] <= 15;
      opCodes[1767] <= 15;
      opCodes[1784] <= 15;
      opCodes[1789] <= 15;
      opCodes[1795] <= 15;
      opCodes[1808] <= 15;
      opCodes[1825] <= 15;
      opCodes[1830] <= 15;
      opCodes[1836] <= 15;
      opCodes[1849] <= 15;
      opCodes[1866] <= 15;
      opCodes[1871] <= 15;
      opCodes[1877] <= 15;
      opCodes[1882] <= 15;
      opCodes[1895] <= 15;
      opCodes[1901] <= 15;
      opCodes[2036] <= 15;
      opCodes[2039] <= 15;
      opCodes[2047] <= 15;
      opCodes[2069] <= 15;
      opCodes[2077] <= 15;
      opCodes[2080] <= 15;
      opCodes[2088] <= 15;
      opCodes[2110] <= 15;
      opCodes[2158] <= 15;
      opCodes[2171] <= 15;
      opCodes[2193] <= 15;
      opCodes[2198] <= 15;
      opCodes[2201] <= 15;
      opCodes[2224] <= 15;
      opCodes[2227] <= 15;
      opCodes[2235] <= 15;
      opCodes[2257] <= 15;
      opCodes[2265] <= 15;
      opCodes[2268] <= 15;
      opCodes[2276] <= 15;
      opCodes[2298] <= 15;
      opCodes[2306] <= 15;
      opCodes[2309] <= 15;
      opCodes[2317] <= 15;
      opCodes[2339] <= 15;
      opCodes[2365] <= 15;
      opCodes[2391] <= 15;
      opCodes[2474] <= 15;
      opCodes[2491] <= 15;
      opCodes[2496] <= 15;
      opCodes[2502] <= 15;
      opCodes[2515] <= 15;
      opCodes[2532] <= 15;
      opCodes[2537] <= 15;
      opCodes[2543] <= 15;
      opCodes[2578] <= 15;
      opCodes[2609] <= 15;
      opCodes[2627] <= 15;
      opCodes[2644] <= 15;
      opCodes[2649] <= 15;
      opCodes[2655] <= 15;
      opCodes[2668] <= 15;
      opCodes[2685] <= 15;
      opCodes[2690] <= 15;
      opCodes[2696] <= 15;
      opCodes[2709] <= 15;
      opCodes[2726] <= 15;
      opCodes[2731] <= 15;
      opCodes[2737] <= 15;
      opCodes[2785] <= 15;
      opCodes[2793] <= 15;
      opCodes[2819] <= 15;
      opCodes[2833] <= 15;
      opCodes[2918] <= 15;
      opCodes[2935] <= 15;
      opCodes[2940] <= 15;
      opCodes[2946] <= 15;
      opCodes[2956] <= 15;
      opCodes[2973] <= 15;
      opCodes[2982] <= 15;
      opCodes[2988] <= 15;
      opCodes[3001] <= 15;
      opCodes[3025] <= 15;
      opCodes[3034] <= 15;
      opCodes[16] <= 16;
      opCodes[54] <= 16;
      opCodes[57] <= 16;
      opCodes[93] <= 16;
      opCodes[174] <= 16;
      opCodes[686] <= 16;
      opCodes[724] <= 16;
      opCodes[727] <= 16;
      opCodes[763] <= 16;
      opCodes[844] <= 16;
      opCodes[913] <= 16;
      opCodes[916] <= 16;
      opCodes[1088] <= 16;
      opCodes[1126] <= 16;
      opCodes[1129] <= 16;
      opCodes[1165] <= 16;
      opCodes[1246] <= 16;
      opCodes[2834] <= 16;
      opCodes[2837] <= 16;
      opCodes[3035] <= 16;
      opCodes[3038] <= 16;
      opCodes[17] <= 17;
      opCodes[30] <= 17;
      opCodes[58] <= 17;
      opCodes[71] <= 17;
      opCodes[94] <= 17;
      opCodes[107] <= 17;
      opCodes[175] <= 17;
      opCodes[188] <= 17;
      opCodes[687] <= 17;
      opCodes[700] <= 17;
      opCodes[728] <= 17;
      opCodes[741] <= 17;
      opCodes[764] <= 17;
      opCodes[777] <= 17;
      opCodes[845] <= 17;
      opCodes[858] <= 17;
      opCodes[917] <= 17;
      opCodes[930] <= 17;
      opCodes[1089] <= 17;
      opCodes[1102] <= 17;
      opCodes[1130] <= 17;
      opCodes[1143] <= 17;
      opCodes[1166] <= 17;
      opCodes[1179] <= 17;
      opCodes[1247] <= 17;
      opCodes[1260] <= 17;
      opCodes[2838] <= 17;
      opCodes[2851] <= 17;
      opCodes[3039] <= 17;
      opCodes[3052] <= 17;
      opCodes[18] <= 18;
      opCodes[31] <= 18;
      opCodes[19] <= 19;
      opCodes[60] <= 19;
      opCodes[96] <= 19;
      opCodes[177] <= 19;
      opCodes[689] <= 19;
      opCodes[730] <= 19;
      opCodes[766] <= 19;
      opCodes[847] <= 19;
      opCodes[919] <= 19;
      opCodes[1091] <= 19;
      opCodes[1132] <= 19;
      opCodes[1168] <= 19;
      opCodes[1249] <= 19;
      opCodes[2840] <= 19;
      opCodes[3041] <= 19;
      opCodes[20] <= 20;
      opCodes[21] <= 21;
      opCodes[62] <= 21;
      opCodes[98] <= 21;
      opCodes[179] <= 21;
      opCodes[691] <= 21;
      opCodes[732] <= 21;
      opCodes[768] <= 21;
      opCodes[849] <= 21;
      opCodes[921] <= 21;
      opCodes[1093] <= 21;
      opCodes[1134] <= 21;
      opCodes[1170] <= 21;
      opCodes[1251] <= 21;
      opCodes[2842] <= 21;
      opCodes[3043] <= 21;
      opCodes[22] <= 22;
      opCodes[63] <= 22;
      opCodes[74] <= 22;
      opCodes[99] <= 22;
      opCodes[180] <= 22;
      opCodes[313] <= 22;
      opCodes[351] <= 22;
      opCodes[387] <= 22;
      opCodes[400] <= 22;
      opCodes[490] <= 22;
      opCodes[528] <= 22;
      opCodes[570] <= 22;
      opCodes[608] <= 22;
      opCodes[692] <= 22;
      opCodes[733] <= 22;
      opCodes[744] <= 22;
      opCodes[769] <= 22;
      opCodes[850] <= 22;
      opCodes[922] <= 22;
      opCodes[933] <= 22;
      opCodes[975] <= 22;
      opCodes[1013] <= 22;
      opCodes[1026] <= 22;
      opCodes[1094] <= 22;
      opCodes[1135] <= 22;
      opCodes[1146] <= 22;
      opCodes[1171] <= 22;
      opCodes[1252] <= 22;
      opCodes[1322] <= 22;
      opCodes[1333] <= 22;
      opCodes[1377] <= 22;
      opCodes[1418] <= 22;
      opCodes[1459] <= 22;
      opCodes[1500] <= 22;
      opCodes[1603] <= 22;
      opCodes[1616] <= 22;
      opCodes[1657] <= 22;
      opCodes[1698] <= 22;
      opCodes[1740] <= 22;
      opCodes[1763] <= 22;
      opCodes[1804] <= 22;
      opCodes[1845] <= 22;
      opCodes[1887] <= 22;
      opCodes[1986] <= 22;
      opCodes[1994] <= 22;
      opCodes[2041] <= 22;
      opCodes[2082] <= 22;
      opCodes[2150] <= 22;
      opCodes[2163] <= 22;
      opCodes[2203] <= 22;
      opCodes[2229] <= 22;
      opCodes[2270] <= 22;
      opCodes[2311] <= 22;
      opCodes[2374] <= 22;
      opCodes[2416] <= 22;
      opCodes[2427] <= 22;
      opCodes[2470] <= 22;
      opCodes[2511] <= 22;
      opCodes[2583] <= 22;
      opCodes[2593] <= 22;
      opCodes[2623] <= 22;
      opCodes[2664] <= 22;
      opCodes[2705] <= 22;
      opCodes[2763] <= 22;
      opCodes[2771] <= 22;
      opCodes[2802] <= 22;
      opCodes[2843] <= 22;
      opCodes[2854] <= 22;
      opCodes[2914] <= 22;
      opCodes[2952] <= 22;
      opCodes[3044] <= 22;
      opCodes[3055] <= 22;
      opCodes[24] <= 23;
      opCodes[65] <= 23;
      opCodes[76] <= 23;
      opCodes[101] <= 23;
      opCodes[182] <= 23;
      opCodes[315] <= 23;
      opCodes[353] <= 23;
      opCodes[389] <= 23;
      opCodes[402] <= 23;
      opCodes[492] <= 23;
      opCodes[530] <= 23;
      opCodes[572] <= 23;
      opCodes[610] <= 23;
      opCodes[694] <= 23;
      opCodes[735] <= 23;
      opCodes[746] <= 23;
      opCodes[771] <= 23;
      opCodes[852] <= 23;
      opCodes[924] <= 23;
      opCodes[935] <= 23;
      opCodes[977] <= 23;
      opCodes[1015] <= 23;
      opCodes[1028] <= 23;
      opCodes[1096] <= 23;
      opCodes[1137] <= 23;
      opCodes[1148] <= 23;
      opCodes[1173] <= 23;
      opCodes[1254] <= 23;
      opCodes[1324] <= 23;
      opCodes[1335] <= 23;
      opCodes[1379] <= 23;
      opCodes[1420] <= 23;
      opCodes[1461] <= 23;
      opCodes[1502] <= 23;
      opCodes[1605] <= 23;
      opCodes[1618] <= 23;
      opCodes[1659] <= 23;
      opCodes[1700] <= 23;
      opCodes[1742] <= 23;
      opCodes[1765] <= 23;
      opCodes[1806] <= 23;
      opCodes[1847] <= 23;
      opCodes[1889] <= 23;
      opCodes[1988] <= 23;
      opCodes[1996] <= 23;
      opCodes[2043] <= 23;
      opCodes[2084] <= 23;
      opCodes[2152] <= 23;
      opCodes[2165] <= 23;
      opCodes[2205] <= 23;
      opCodes[2231] <= 23;
      opCodes[2272] <= 23;
      opCodes[2313] <= 23;
      opCodes[2376] <= 23;
      opCodes[2418] <= 23;
      opCodes[2429] <= 23;
      opCodes[2472] <= 23;
      opCodes[2513] <= 23;
      opCodes[2585] <= 23;
      opCodes[2595] <= 23;
      opCodes[2625] <= 23;
      opCodes[2666] <= 23;
      opCodes[2707] <= 23;
      opCodes[2765] <= 23;
      opCodes[2773] <= 23;
      opCodes[2804] <= 23;
      opCodes[2845] <= 23;
      opCodes[2856] <= 23;
      opCodes[2916] <= 23;
      opCodes[2954] <= 23;
      opCodes[3046] <= 23;
      opCodes[3057] <= 23;
      opCodes[25] <= 24;
      opCodes[66] <= 24;
      opCodes[77] <= 24;
      opCodes[102] <= 24;
      opCodes[140] <= 24;
      opCodes[183] <= 24;
      opCodes[196] <= 24;
      opCodes[316] <= 24;
      opCodes[354] <= 24;
      opCodes[390] <= 24;
      opCodes[403] <= 24;
      opCodes[420] <= 24;
      opCodes[433] <= 24;
      opCodes[493] <= 24;
      opCodes[531] <= 24;
      opCodes[573] <= 24;
      opCodes[611] <= 24;
      opCodes[651] <= 24;
      opCodes[664] <= 24;
      opCodes[695] <= 24;
      opCodes[736] <= 24;
      opCodes[747] <= 24;
      opCodes[772] <= 24;
      opCodes[810] <= 24;
      opCodes[853] <= 24;
      opCodes[866] <= 24;
      opCodes[925] <= 24;
      opCodes[936] <= 24;
      opCodes[978] <= 24;
      opCodes[1016] <= 24;
      opCodes[1029] <= 24;
      opCodes[1044] <= 24;
      opCodes[1097] <= 24;
      opCodes[1138] <= 24;
      opCodes[1149] <= 24;
      opCodes[1174] <= 24;
      opCodes[1212] <= 24;
      opCodes[1255] <= 24;
      opCodes[1268] <= 24;
      opCodes[1325] <= 24;
      opCodes[1336] <= 24;
      opCodes[1380] <= 24;
      opCodes[1421] <= 24;
      opCodes[1462] <= 24;
      opCodes[1503] <= 24;
      opCodes[1606] <= 24;
      opCodes[1619] <= 24;
      opCodes[1660] <= 24;
      opCodes[1701] <= 24;
      opCodes[1743] <= 24;
      opCodes[1766] <= 24;
      opCodes[1807] <= 24;
      opCodes[1848] <= 24;
      opCodes[1890] <= 24;
      opCodes[1989] <= 24;
      opCodes[1997] <= 24;
      opCodes[2044] <= 24;
      opCodes[2085] <= 24;
      opCodes[2153] <= 24;
      opCodes[2166] <= 24;
      opCodes[2206] <= 24;
      opCodes[2232] <= 24;
      opCodes[2273] <= 24;
      opCodes[2314] <= 24;
      opCodes[2377] <= 24;
      opCodes[2419] <= 24;
      opCodes[2430] <= 24;
      opCodes[2473] <= 24;
      opCodes[2514] <= 24;
      opCodes[2586] <= 24;
      opCodes[2596] <= 24;
      opCodes[2600] <= 24;
      opCodes[2626] <= 24;
      opCodes[2667] <= 24;
      opCodes[2708] <= 24;
      opCodes[2766] <= 24;
      opCodes[2774] <= 24;
      opCodes[2805] <= 24;
      opCodes[2846] <= 24;
      opCodes[2857] <= 24;
      opCodes[2917] <= 24;
      opCodes[2955] <= 24;
      opCodes[2996] <= 24;
      opCodes[3047] <= 24;
      opCodes[3058] <= 24;
      opCodes[26] <= 25;
      opCodes[27] <= 26;
      opCodes[37] <= 26;
      opCodes[68] <= 26;
      opCodes[104] <= 26;
      opCodes[116] <= 26;
      opCodes[185] <= 26;
      opCodes[197] <= 26;
      opCodes[397] <= 26;
      opCodes[697] <= 26;
      opCodes[707] <= 26;
      opCodes[738] <= 26;
      opCodes[774] <= 26;
      opCodes[786] <= 26;
      opCodes[855] <= 26;
      opCodes[867] <= 26;
      opCodes[927] <= 26;
      opCodes[949] <= 26;
      opCodes[1023] <= 26;
      opCodes[1047] <= 26;
      opCodes[1099] <= 26;
      opCodes[1109] <= 26;
      opCodes[1140] <= 26;
      opCodes[1176] <= 26;
      opCodes[1188] <= 26;
      opCodes[1257] <= 26;
      opCodes[1269] <= 26;
      opCodes[1330] <= 26;
      opCodes[1737] <= 26;
      opCodes[1884] <= 26;
      opCodes[1983] <= 26;
      opCodes[2147] <= 26;
      opCodes[2160] <= 26;
      opCodes[2362] <= 26;
      opCodes[2367] <= 26;
      opCodes[2424] <= 26;
      opCodes[2580] <= 26;
      opCodes[2760] <= 26;
      opCodes[2790] <= 26;
      opCodes[2795] <= 26;
      opCodes[2848] <= 26;
      opCodes[2888] <= 26;
      opCodes[2999] <= 26;
      opCodes[3049] <= 26;
      opCodes[28] <= 27;
      opCodes[69] <= 27;
      opCodes[105] <= 27;
      opCodes[126] <= 27;
      opCodes[150] <= 27;
      opCodes[186] <= 27;
      opCodes[224] <= 27;
      opCodes[328] <= 27;
      opCodes[331] <= 27;
      opCodes[346] <= 27;
      opCodes[366] <= 27;
      opCodes[369] <= 27;
      opCodes[384] <= 27;
      opCodes[428] <= 27;
      opCodes[441] <= 27;
      opCodes[505] <= 27;
      opCodes[508] <= 27;
      opCodes[523] <= 27;
      opCodes[543] <= 27;
      opCodes[546] <= 27;
      opCodes[565] <= 27;
      opCodes[585] <= 27;
      opCodes[588] <= 27;
      opCodes[603] <= 27;
      opCodes[623] <= 27;
      opCodes[626] <= 27;
      opCodes[643] <= 27;
      opCodes[659] <= 27;
      opCodes[672] <= 27;
      opCodes[698] <= 27;
      opCodes[739] <= 27;
      opCodes[775] <= 27;
      opCodes[796] <= 27;
      opCodes[820] <= 27;
      opCodes[856] <= 27;
      opCodes[894] <= 27;
      opCodes[928] <= 27;
      opCodes[990] <= 27;
      opCodes[993] <= 27;
      opCodes[1008] <= 27;
      opCodes[1074] <= 27;
      opCodes[1100] <= 27;
      opCodes[1141] <= 27;
      opCodes[1177] <= 27;
      opCodes[1198] <= 27;
      opCodes[1222] <= 27;
      opCodes[1258] <= 27;
      opCodes[1296] <= 27;
      opCodes[1392] <= 27;
      opCodes[1395] <= 27;
      opCodes[1410] <= 27;
      opCodes[1433] <= 27;
      opCodes[1436] <= 27;
      opCodes[1451] <= 27;
      opCodes[1474] <= 27;
      opCodes[1477] <= 27;
      opCodes[1492] <= 27;
      opCodes[1515] <= 27;
      opCodes[1518] <= 27;
      opCodes[1533] <= 27;
      opCodes[1595] <= 27;
      opCodes[1631] <= 27;
      opCodes[1634] <= 27;
      opCodes[1649] <= 27;
      opCodes[1672] <= 27;
      opCodes[1675] <= 27;
      opCodes[1690] <= 27;
      opCodes[1713] <= 27;
      opCodes[1716] <= 27;
      opCodes[1731] <= 27;
      opCodes[1755] <= 27;
      opCodes[1778] <= 27;
      opCodes[1781] <= 27;
      opCodes[1796] <= 27;
      opCodes[1819] <= 27;
      opCodes[1822] <= 27;
      opCodes[1837] <= 27;
      opCodes[1860] <= 27;
      opCodes[1863] <= 27;
      opCodes[1878] <= 27;
      opCodes[1902] <= 27;
      opCodes[1956] <= 27;
      opCodes[2070] <= 27;
      opCodes[2111] <= 27;
      opCodes[2136] <= 27;
      opCodes[2194] <= 27;
      opCodes[2217] <= 27;
      opCodes[2258] <= 27;
      opCodes[2299] <= 27;
      opCodes[2340] <= 27;
      opCodes[2372] <= 27;
      opCodes[2385] <= 27;
      opCodes[2388] <= 27;
      opCodes[2425] <= 27;
      opCodes[2485] <= 27;
      opCodes[2488] <= 27;
      opCodes[2503] <= 27;
      opCodes[2526] <= 27;
      opCodes[2529] <= 27;
      opCodes[2544] <= 27;
      opCodes[2569] <= 27;
      opCodes[2610] <= 27;
      opCodes[2615] <= 27;
      opCodes[2638] <= 27;
      opCodes[2641] <= 27;
      opCodes[2656] <= 27;
      opCodes[2679] <= 27;
      opCodes[2682] <= 27;
      opCodes[2697] <= 27;
      opCodes[2720] <= 27;
      opCodes[2723] <= 27;
      opCodes[2738] <= 27;
      opCodes[2761] <= 27;
      opCodes[2786] <= 27;
      opCodes[2791] <= 27;
      opCodes[2800] <= 27;
      opCodes[2813] <= 27;
      opCodes[2816] <= 27;
      opCodes[2824] <= 27;
      opCodes[2849] <= 27;
      opCodes[2861] <= 27;
      opCodes[2929] <= 27;
      opCodes[2932] <= 27;
      opCodes[2947] <= 27;
      opCodes[2967] <= 27;
      opCodes[2970] <= 27;
      opCodes[2989] <= 27;
      opCodes[3026] <= 27;
      opCodes[3050] <= 27;
      opCodes[3066] <= 27;
      opCodes[29] <= 28;
      opCodes[70] <= 28;
      opCodes[106] <= 28;
      opCodes[142] <= 28;
      opCodes[187] <= 28;
      opCodes[340] <= 28;
      opCodes[378] <= 28;
      opCodes[396] <= 28;
      opCodes[399] <= 28;
      opCodes[422] <= 28;
      opCodes[435] <= 28;
      opCodes[517] <= 28;
      opCodes[559] <= 28;
      opCodes[597] <= 28;
      opCodes[637] <= 28;
      opCodes[653] <= 28;
      opCodes[666] <= 28;
      opCodes[699] <= 28;
      opCodes[740] <= 28;
      opCodes[776] <= 28;
      opCodes[812] <= 28;
      opCodes[857] <= 28;
      opCodes[929] <= 28;
      opCodes[1002] <= 28;
      opCodes[1022] <= 28;
      opCodes[1025] <= 28;
      opCodes[1046] <= 28;
      opCodes[1101] <= 28;
      opCodes[1142] <= 28;
      opCodes[1178] <= 28;
      opCodes[1214] <= 28;
      opCodes[1259] <= 28;
      opCodes[1329] <= 28;
      opCodes[1332] <= 28;
      opCodes[1404] <= 28;
      opCodes[1445] <= 28;
      opCodes[1486] <= 28;
      opCodes[1527] <= 28;
      opCodes[1643] <= 28;
      opCodes[1684] <= 28;
      opCodes[1725] <= 28;
      opCodes[1736] <= 28;
      opCodes[1739] <= 28;
      opCodes[1749] <= 28;
      opCodes[1790] <= 28;
      opCodes[1831] <= 28;
      opCodes[1872] <= 28;
      opCodes[1883] <= 28;
      opCodes[1886] <= 28;
      opCodes[1896] <= 28;
      opCodes[1982] <= 28;
      opCodes[1985] <= 28;
      opCodes[1993] <= 28;
      opCodes[2040] <= 28;
      opCodes[2081] <= 28;
      opCodes[2146] <= 28;
      opCodes[2149] <= 28;
      opCodes[2159] <= 28;
      opCodes[2162] <= 28;
      opCodes[2202] <= 28;
      opCodes[2228] <= 28;
      opCodes[2269] <= 28;
      opCodes[2310] <= 28;
      opCodes[2361] <= 28;
      opCodes[2364] <= 28;
      opCodes[2415] <= 28;
      opCodes[2423] <= 28;
      opCodes[2426] <= 28;
      opCodes[2497] <= 28;
      opCodes[2538] <= 28;
      opCodes[2579] <= 28;
      opCodes[2582] <= 28;
      opCodes[2592] <= 28;
      opCodes[2602] <= 28;
      opCodes[2650] <= 28;
      opCodes[2691] <= 28;
      opCodes[2732] <= 28;
      opCodes[2759] <= 28;
      opCodes[2762] <= 28;
      opCodes[2770] <= 28;
      opCodes[2778] <= 28;
      opCodes[2789] <= 28;
      opCodes[2792] <= 28;
      opCodes[2850] <= 28;
      opCodes[2941] <= 28;
      opCodes[2983] <= 28;
      opCodes[2998] <= 28;
      opCodes[3051] <= 28;
      opCodes[32] <= 29;
      opCodes[33] <= 30;
      opCodes[44] <= 30;
      opCodes[310] <= 30;
      opCodes[348] <= 30;
      opCodes[414] <= 30;
      opCodes[430] <= 30;
      opCodes[487] <= 30;
      opCodes[525] <= 30;
      opCodes[556] <= 30;
      opCodes[567] <= 30;
      opCodes[605] <= 30;
      opCodes[634] <= 30;
      opCodes[645] <= 30;
      opCodes[661] <= 30;
      opCodes[703] <= 30;
      opCodes[714] <= 30;
      opCodes[903] <= 30;
      opCodes[1105] <= 30;
      opCodes[1116] <= 30;
      opCodes[1339] <= 30;
      opCodes[1368] <= 30;
      opCodes[1401] <= 30;
      opCodes[1442] <= 30;
      opCodes[1483] <= 30;
      opCodes[1524] <= 30;
      opCodes[1535] <= 30;
      opCodes[1600] <= 30;
      opCodes[1640] <= 30;
      opCodes[1681] <= 30;
      opCodes[1722] <= 30;
      opCodes[1744] <= 30;
      opCodes[1787] <= 30;
      opCodes[1828] <= 30;
      opCodes[1869] <= 30;
      opCodes[1891] <= 30;
      opCodes[1893] <= 30;
      opCodes[1936] <= 30;
      opCodes[2980] <= 30;
      opCodes[34] <= 31;
      opCodes[113] <= 31;
      opCodes[704] <= 31;
      opCodes[783] <= 31;
      opCodes[1106] <= 31;
      opCodes[1185] <= 31;
      opCodes[35] <= 32;
      opCodes[114] <= 32;
      opCodes[705] <= 32;
      opCodes[784] <= 32;
      opCodes[1107] <= 32;
      opCodes[1186] <= 32;
      opCodes[36] <= 33;
      opCodes[115] <= 33;
      opCodes[706] <= 33;
      opCodes[785] <= 33;
      opCodes[1108] <= 33;
      opCodes[1187] <= 33;
      opCodes[38] <= 34;
      opCodes[117] <= 34;
      opCodes[708] <= 34;
      opCodes[787] <= 34;
      opCodes[1110] <= 34;
      opCodes[1189] <= 34;
      opCodes[39] <= 35;
      opCodes[118] <= 35;
      opCodes[143] <= 35;
      opCodes[219] <= 35;
      opCodes[341] <= 35;
      opCodes[379] <= 35;
      opCodes[391] <= 35;
      opCodes[404] <= 35;
      opCodes[423] <= 35;
      opCodes[436] <= 35;
      opCodes[518] <= 35;
      opCodes[552] <= 35;
      opCodes[560] <= 35;
      opCodes[598] <= 35;
      opCodes[638] <= 35;
      opCodes[654] <= 35;
      opCodes[667] <= 35;
      opCodes[709] <= 35;
      opCodes[788] <= 35;
      opCodes[813] <= 35;
      opCodes[889] <= 35;
      opCodes[1003] <= 35;
      opCodes[1017] <= 35;
      opCodes[1030] <= 35;
      opCodes[1069] <= 35;
      opCodes[1111] <= 35;
      opCodes[1190] <= 35;
      opCodes[1215] <= 35;
      opCodes[1291] <= 35;
      opCodes[1405] <= 35;
      opCodes[1446] <= 35;
      opCodes[1487] <= 35;
      opCodes[1528] <= 35;
      opCodes[1607] <= 35;
      opCodes[1644] <= 35;
      opCodes[1685] <= 35;
      opCodes[1726] <= 35;
      opCodes[1750] <= 35;
      opCodes[1791] <= 35;
      opCodes[1832] <= 35;
      opCodes[1873] <= 35;
      opCodes[1897] <= 35;
      opCodes[2065] <= 35;
      opCodes[2106] <= 35;
      opCodes[2154] <= 35;
      opCodes[2189] <= 35;
      opCodes[2253] <= 35;
      opCodes[2294] <= 35;
      opCodes[2335] <= 35;
      opCodes[2498] <= 35;
      opCodes[2539] <= 35;
      opCodes[2603] <= 35;
      opCodes[2651] <= 35;
      opCodes[2692] <= 35;
      opCodes[2733] <= 35;
      opCodes[2767] <= 35;
      opCodes[2779] <= 35;
      opCodes[2942] <= 35;
      opCodes[2976] <= 35;
      opCodes[2984] <= 35;
      opCodes[3021] <= 35;
      opCodes[40] <= 36;
      opCodes[119] <= 36;
      opCodes[710] <= 36;
      opCodes[789] <= 36;
      opCodes[1112] <= 36;
      opCodes[1191] <= 36;
      opCodes[41] <= 37;
      opCodes[78] <= 37;
      opCodes[120] <= 37;
      opCodes[145] <= 37;
      opCodes[221] <= 37;
      opCodes[343] <= 37;
      opCodes[381] <= 37;
      opCodes[425] <= 37;
      opCodes[438] <= 37;
      opCodes[520] <= 37;
      opCodes[562] <= 37;
      opCodes[600] <= 37;
      opCodes[640] <= 37;
      opCodes[656] <= 37;
      opCodes[669] <= 37;
      opCodes[711] <= 37;
      opCodes[748] <= 37;
      opCodes[790] <= 37;
      opCodes[815] <= 37;
      opCodes[891] <= 37;
      opCodes[937] <= 37;
      opCodes[1005] <= 37;
      opCodes[1071] <= 37;
      opCodes[1113] <= 37;
      opCodes[1150] <= 37;
      opCodes[1192] <= 37;
      opCodes[1217] <= 37;
      opCodes[1293] <= 37;
      opCodes[1326] <= 37;
      opCodes[1337] <= 37;
      opCodes[1407] <= 37;
      opCodes[1448] <= 37;
      opCodes[1489] <= 37;
      opCodes[1530] <= 37;
      opCodes[1646] <= 37;
      opCodes[1687] <= 37;
      opCodes[1728] <= 37;
      opCodes[1752] <= 37;
      opCodes[1793] <= 37;
      opCodes[1834] <= 37;
      opCodes[1875] <= 37;
      opCodes[1899] <= 37;
      opCodes[1990] <= 37;
      opCodes[1998] <= 37;
      opCodes[2067] <= 37;
      opCodes[2108] <= 37;
      opCodes[2191] <= 37;
      opCodes[2255] <= 37;
      opCodes[2296] <= 37;
      opCodes[2337] <= 37;
      opCodes[2420] <= 37;
      opCodes[2431] <= 37;
      opCodes[2500] <= 37;
      opCodes[2541] <= 37;
      opCodes[2587] <= 37;
      opCodes[2605] <= 37;
      opCodes[2653] <= 37;
      opCodes[2694] <= 37;
      opCodes[2735] <= 37;
      opCodes[2781] <= 37;
      opCodes[2858] <= 37;
      opCodes[2944] <= 37;
      opCodes[2986] <= 37;
      opCodes[3023] <= 37;
      opCodes[3059] <= 37;
      opCodes[42] <= 38;
      opCodes[121] <= 38;
      opCodes[712] <= 38;
      opCodes[791] <= 38;
      opCodes[1114] <= 38;
      opCodes[1193] <= 38;
      opCodes[43] <= 39;
      opCodes[122] <= 39;
      opCodes[45] <= 40;
      opCodes[124] <= 40;
      opCodes[715] <= 40;
      opCodes[794] <= 40;
      opCodes[904] <= 40;
      opCodes[1117] <= 40;
      opCodes[1196] <= 40;
      opCodes[1937] <= 40;
      opCodes[2859] <= 40;
      opCodes[3060] <= 40;
      opCodes[3064] <= 40;
      opCodes[46] <= 41;
      opCodes[716] <= 41;
      opCodes[1118] <= 41;
      opCodes[47] <= 42;
      opCodes[717] <= 42;
      opCodes[906] <= 42;
      opCodes[947] <= 42;
      opCodes[1119] <= 42;
      opCodes[1940] <= 42;
      opCodes[1946] <= 42;
      opCodes[1961] <= 42;
      opCodes[2400] <= 42;
      opCodes[2827] <= 42;
      opCodes[2886] <= 42;
      opCodes[3028] <= 42;
      opCodes[48] <= 43;
      opCodes[87] <= 43;
      opCodes[136] <= 43;
      opCodes[168] <= 43;
      opCodes[192] <= 43;
      opCodes[311] <= 43;
      opCodes[338] <= 43;
      opCodes[349] <= 43;
      opCodes[376] <= 43;
      opCodes[394] <= 43;
      opCodes[415] <= 43;
      opCodes[488] <= 43;
      opCodes[515] <= 43;
      opCodes[526] <= 43;
      opCodes[555] <= 43;
      opCodes[568] <= 43;
      opCodes[595] <= 43;
      opCodes[606] <= 43;
      opCodes[633] <= 43;
      opCodes[646] <= 43;
      opCodes[718] <= 43;
      opCodes[757] <= 43;
      opCodes[806] <= 43;
      opCodes[838] <= 43;
      opCodes[862] <= 43;
      opCodes[907] <= 43;
      opCodes[973] <= 43;
      opCodes[1000] <= 43;
      opCodes[1011] <= 43;
      opCodes[1020] <= 43;
      opCodes[1040] <= 43;
      opCodes[1120] <= 43;
      opCodes[1159] <= 43;
      opCodes[1208] <= 43;
      opCodes[1240] <= 43;
      opCodes[1264] <= 43;
      opCodes[1369] <= 43;
      opCodes[1375] <= 43;
      opCodes[1402] <= 43;
      opCodes[1416] <= 43;
      opCodes[1443] <= 43;
      opCodes[1457] <= 43;
      opCodes[1484] <= 43;
      opCodes[1498] <= 43;
      opCodes[1525] <= 43;
      opCodes[1601] <= 43;
      opCodes[1614] <= 43;
      opCodes[1641] <= 43;
      opCodes[1655] <= 43;
      opCodes[1682] <= 43;
      opCodes[1696] <= 43;
      opCodes[1723] <= 43;
      opCodes[1734] <= 43;
      opCodes[1745] <= 43;
      opCodes[1761] <= 43;
      opCodes[1788] <= 43;
      opCodes[1802] <= 43;
      opCodes[1829] <= 43;
      opCodes[1843] <= 43;
      opCodes[1870] <= 43;
      opCodes[1881] <= 43;
      opCodes[1892] <= 43;
      opCodes[1980] <= 43;
      opCodes[2035] <= 43;
      opCodes[2046] <= 43;
      opCodes[2076] <= 43;
      opCodes[2087] <= 43;
      opCodes[2144] <= 43;
      opCodes[2157] <= 43;
      opCodes[2168] <= 43;
      opCodes[2197] <= 43;
      opCodes[2223] <= 43;
      opCodes[2234] <= 43;
      opCodes[2264] <= 43;
      opCodes[2275] <= 43;
      opCodes[2305] <= 43;
      opCodes[2316] <= 43;
      opCodes[2359] <= 43;
      opCodes[2413] <= 43;
      opCodes[2468] <= 43;
      opCodes[2495] <= 43;
      opCodes[2509] <= 43;
      opCodes[2536] <= 43;
      opCodes[2577] <= 43;
      opCodes[2590] <= 43;
      opCodes[2598] <= 43;
      opCodes[2621] <= 43;
      opCodes[2648] <= 43;
      opCodes[2662] <= 43;
      opCodes[2689] <= 43;
      opCodes[2703] <= 43;
      opCodes[2730] <= 43;
      opCodes[2757] <= 43;
      opCodes[2828] <= 43;
      opCodes[2912] <= 43;
      opCodes[2939] <= 43;
      opCodes[2950] <= 43;
      opCodes[2979] <= 43;
      opCodes[2992] <= 43;
      opCodes[3029] <= 43;
      opCodes[55] <= 44;
      opCodes[725] <= 44;
      opCodes[914] <= 44;
      opCodes[1127] <= 44;
      opCodes[2835] <= 44;
      opCodes[3036] <= 44;
      opCodes[56] <= 45;
      opCodes[204] <= 45;
      opCodes[213] <= 45;
      opCodes[216] <= 45;
      opCodes[254] <= 45;
      opCodes[335] <= 45;
      opCodes[373] <= 45;
      opCodes[398] <= 45;
      opCodes[512] <= 45;
      opCodes[550] <= 45;
      opCodes[592] <= 45;
      opCodes[630] <= 45;
      opCodes[726] <= 45;
      opCodes[874] <= 45;
      opCodes[883] <= 45;
      opCodes[886] <= 45;
      opCodes[915] <= 45;
      opCodes[997] <= 45;
      opCodes[1024] <= 45;
      opCodes[1054] <= 45;
      opCodes[1063] <= 45;
      opCodes[1066] <= 45;
      opCodes[1128] <= 45;
      opCodes[1276] <= 45;
      opCodes[1285] <= 45;
      opCodes[1288] <= 45;
      opCodes[1313] <= 45;
      opCodes[1331] <= 45;
      opCodes[1399] <= 45;
      opCodes[1440] <= 45;
      opCodes[1481] <= 45;
      opCodes[1522] <= 45;
      opCodes[1577] <= 45;
      opCodes[1586] <= 45;
      opCodes[1638] <= 45;
      opCodes[1679] <= 45;
      opCodes[1720] <= 45;
      opCodes[1738] <= 45;
      opCodes[1785] <= 45;
      opCodes[1826] <= 45;
      opCodes[1867] <= 45;
      opCodes[1885] <= 45;
      opCodes[1951] <= 45;
      opCodes[1973] <= 45;
      opCodes[1984] <= 45;
      opCodes[2037] <= 45;
      opCodes[2054] <= 45;
      opCodes[2061] <= 45;
      opCodes[2078] <= 45;
      opCodes[2095] <= 45;
      opCodes[2102] <= 45;
      opCodes[2120] <= 45;
      opCodes[2129] <= 45;
      opCodes[2148] <= 45;
      opCodes[2161] <= 45;
      opCodes[2178] <= 45;
      opCodes[2185] <= 45;
      opCodes[2199] <= 45;
      opCodes[2212] <= 45;
      opCodes[2225] <= 45;
      opCodes[2242] <= 45;
      opCodes[2249] <= 45;
      opCodes[2266] <= 45;
      opCodes[2283] <= 45;
      opCodes[2290] <= 45;
      opCodes[2307] <= 45;
      opCodes[2324] <= 45;
      opCodes[2331] <= 45;
      opCodes[2363] <= 45;
      opCodes[2392] <= 45;
      opCodes[2398] <= 45;
      opCodes[2408] <= 45;
      opCodes[2492] <= 45;
      opCodes[2533] <= 45;
      opCodes[2553] <= 45;
      opCodes[2562] <= 45;
      opCodes[2581] <= 45;
      opCodes[2645] <= 45;
      opCodes[2686] <= 45;
      opCodes[2727] <= 45;
      opCodes[2820] <= 45;
      opCodes[2836] <= 45;
      opCodes[2876] <= 45;
      opCodes[2936] <= 45;
      opCodes[2974] <= 45;
      opCodes[3006] <= 45;
      opCodes[3015] <= 45;
      opCodes[3018] <= 45;
      opCodes[3037] <= 45;
      opCodes[59] <= 46;
      opCodes[72] <= 46;
      opCodes[61] <= 47;
      opCodes[67] <= 48;
      opCodes[73] <= 49;
      opCodes[79] <= 50;
      opCodes[749] <= 50;
      opCodes[938] <= 50;
      opCodes[1151] <= 50;
      opCodes[80] <= 51;
      opCodes[86] <= 51;
      opCodes[110] <= 51;
      opCodes[123] <= 51;
      opCodes[750] <= 51;
      opCodes[756] <= 51;
      opCodes[780] <= 51;
      opCodes[793] <= 51;
      opCodes[939] <= 51;
      opCodes[945] <= 51;
      opCodes[1152] <= 51;
      opCodes[1158] <= 51;
      opCodes[1182] <= 51;
      opCodes[1195] <= 51;
      opCodes[2869] <= 51;
      opCodes[2884] <= 51;
      opCodes[3063] <= 51;
      opCodes[81] <= 52;
      opCodes[83] <= 52;
      opCodes[235] <= 52;
      opCodes[237] <= 52;
      opCodes[751] <= 52;
      opCodes[753] <= 52;
      opCodes[940] <= 52;
      opCodes[942] <= 52;
      opCodes[1153] <= 52;
      opCodes[1155] <= 52;
      opCodes[1342] <= 52;
      opCodes[1344] <= 52;
      opCodes[1941] <= 52;
      opCodes[1943] <= 52;
      opCodes[2003] <= 52;
      opCodes[2005] <= 52;
      opCodes[2436] <= 52;
      opCodes[2438] <= 52;
      opCodes[82] <= 53;
      opCodes[236] <= 53;
      opCodes[752] <= 53;
      opCodes[941] <= 53;
      opCodes[1154] <= 53;
      opCodes[1343] <= 53;
      opCodes[1942] <= 53;
      opCodes[2004] <= 53;
      opCodes[2437] <= 53;
      opCodes[84] <= 54;
      opCodes[238] <= 54;
      opCodes[754] <= 54;
      opCodes[943] <= 54;
      opCodes[1156] <= 54;
      opCodes[1345] <= 54;
      opCodes[1944] <= 54;
      opCodes[2006] <= 54;
      opCodes[2439] <= 54;
      opCodes[85] <= 55;
      opCodes[95] <= 56;
      opCodes[108] <= 56;
      opCodes[97] <= 57;
      opCodes[103] <= 58;
      opCodes[109] <= 59;
      opCodes[111] <= 60;
      opCodes[781] <= 60;
      opCodes[1183] <= 60;
      opCodes[112] <= 61;
      opCodes[782] <= 61;
      opCodes[1184] <= 61;
      opCodes[125] <= 62;
      opCodes[128] <= 62;
      opCodes[795] <= 62;
      opCodes[798] <= 62;
      opCodes[1197] <= 62;
      opCodes[1200] <= 62;
      opCodes[127] <= 63;
      opCodes[797] <= 63;
      opCodes[1199] <= 63;
      opCodes[129] <= 64;
      opCodes[799] <= 64;
      opCodes[1201] <= 64;
      opCodes[2864] <= 64;
      opCodes[3069] <= 64;
      opCodes[130] <= 65;
      opCodes[131] <= 66;
      opCodes[132] <= 67;
      opCodes[272] <= 67;
      opCodes[293] <= 67;
      opCodes[449] <= 67;
      opCodes[470] <= 67;
      opCodes[802] <= 67;
      opCodes[955] <= 67;
      opCodes[1204] <= 67;
      opCodes[2867] <= 67;
      opCodes[2894] <= 67;
      opCodes[3072] <= 67;
      opCodes[133] <= 68;
      opCodes[803] <= 68;
      opCodes[1205] <= 68;
      opCodes[134] <= 69;
      opCodes[135] <= 70;
      opCodes[155] <= 70;
      opCodes[167] <= 70;
      opCodes[191] <= 70;
      opCodes[805] <= 70;
      opCodes[825] <= 70;
      opCodes[837] <= 70;
      opCodes[861] <= 70;
      opCodes[1207] <= 70;
      opCodes[1227] <= 70;
      opCodes[1239] <= 70;
      opCodes[1263] <= 70;
      opCodes[139] <= 71;
      opCodes[195] <= 71;
      opCodes[809] <= 71;
      opCodes[865] <= 71;
      opCodes[1211] <= 71;
      opCodes[1267] <= 71;
      opCodes[141] <= 72;
      opCodes[811] <= 72;
      opCodes[1213] <= 72;
      opCodes[144] <= 73;
      opCodes[220] <= 73;
      opCodes[342] <= 73;
      opCodes[380] <= 73;
      opCodes[424] <= 73;
      opCodes[437] <= 73;
      opCodes[519] <= 73;
      opCodes[561] <= 73;
      opCodes[599] <= 73;
      opCodes[639] <= 73;
      opCodes[655] <= 73;
      opCodes[668] <= 73;
      opCodes[814] <= 73;
      opCodes[890] <= 73;
      opCodes[1004] <= 73;
      opCodes[1070] <= 73;
      opCodes[1216] <= 73;
      opCodes[1292] <= 73;
      opCodes[1406] <= 73;
      opCodes[1447] <= 73;
      opCodes[1488] <= 73;
      opCodes[1529] <= 73;
      opCodes[1645] <= 73;
      opCodes[1686] <= 73;
      opCodes[1727] <= 73;
      opCodes[1751] <= 73;
      opCodes[1792] <= 73;
      opCodes[1833] <= 73;
      opCodes[1874] <= 73;
      opCodes[1898] <= 73;
      opCodes[2066] <= 73;
      opCodes[2107] <= 73;
      opCodes[2190] <= 73;
      opCodes[2254] <= 73;
      opCodes[2295] <= 73;
      opCodes[2336] <= 73;
      opCodes[2499] <= 73;
      opCodes[2540] <= 73;
      opCodes[2604] <= 73;
      opCodes[2652] <= 73;
      opCodes[2693] <= 73;
      opCodes[2734] <= 73;
      opCodes[2780] <= 73;
      opCodes[2943] <= 73;
      opCodes[2985] <= 73;
      opCodes[3022] <= 73;
      opCodes[146] <= 74;
      opCodes[222] <= 74;
      opCodes[344] <= 74;
      opCodes[382] <= 74;
      opCodes[426] <= 74;
      opCodes[439] <= 74;
      opCodes[521] <= 74;
      opCodes[563] <= 74;
      opCodes[601] <= 74;
      opCodes[641] <= 74;
      opCodes[657] <= 74;
      opCodes[670] <= 74;
      opCodes[816] <= 74;
      opCodes[892] <= 74;
      opCodes[1006] <= 74;
      opCodes[1072] <= 74;
      opCodes[1218] <= 74;
      opCodes[1294] <= 74;
      opCodes[1408] <= 74;
      opCodes[1449] <= 74;
      opCodes[1490] <= 74;
      opCodes[1531] <= 74;
      opCodes[1647] <= 74;
      opCodes[1688] <= 74;
      opCodes[1729] <= 74;
      opCodes[1753] <= 74;
      opCodes[1794] <= 74;
      opCodes[1835] <= 74;
      opCodes[1876] <= 74;
      opCodes[1900] <= 74;
      opCodes[2068] <= 74;
      opCodes[2109] <= 74;
      opCodes[2192] <= 74;
      opCodes[2256] <= 74;
      opCodes[2297] <= 74;
      opCodes[2338] <= 74;
      opCodes[2501] <= 74;
      opCodes[2542] <= 74;
      opCodes[2606] <= 74;
      opCodes[2654] <= 74;
      opCodes[2695] <= 74;
      opCodes[2736] <= 74;
      opCodes[2782] <= 74;
      opCodes[2945] <= 74;
      opCodes[2987] <= 74;
      opCodes[3024] <= 74;
      opCodes[147] <= 75;
      opCodes[817] <= 75;
      opCodes[1219] <= 75;
      opCodes[2607] <= 75;
      opCodes[2783] <= 75;
      opCodes[148] <= 76;
      opCodes[151] <= 77;
      opCodes[225] <= 77;
      opCodes[336] <= 77;
      opCodes[347] <= 77;
      opCodes[374] <= 77;
      opCodes[385] <= 77;
      opCodes[429] <= 77;
      opCodes[442] <= 77;
      opCodes[513] <= 77;
      opCodes[524] <= 77;
      opCodes[551] <= 77;
      opCodes[566] <= 77;
      opCodes[593] <= 77;
      opCodes[604] <= 77;
      opCodes[631] <= 77;
      opCodes[644] <= 77;
      opCodes[660] <= 77;
      opCodes[673] <= 77;
      opCodes[821] <= 77;
      opCodes[895] <= 77;
      opCodes[998] <= 77;
      opCodes[1009] <= 77;
      opCodes[1075] <= 77;
      opCodes[1223] <= 77;
      opCodes[1297] <= 77;
      opCodes[1400] <= 77;
      opCodes[1411] <= 77;
      opCodes[1441] <= 77;
      opCodes[1452] <= 77;
      opCodes[1482] <= 77;
      opCodes[1493] <= 77;
      opCodes[1523] <= 77;
      opCodes[1534] <= 77;
      opCodes[1639] <= 77;
      opCodes[1650] <= 77;
      opCodes[1680] <= 77;
      opCodes[1691] <= 77;
      opCodes[1721] <= 77;
      opCodes[1732] <= 77;
      opCodes[1756] <= 77;
      opCodes[1786] <= 77;
      opCodes[1797] <= 77;
      opCodes[1827] <= 77;
      opCodes[1838] <= 77;
      opCodes[1868] <= 77;
      opCodes[1879] <= 77;
      opCodes[1903] <= 77;
      opCodes[2038] <= 77;
      opCodes[2071] <= 77;
      opCodes[2079] <= 77;
      opCodes[2112] <= 77;
      opCodes[2195] <= 77;
      opCodes[2200] <= 77;
      opCodes[2226] <= 77;
      opCodes[2259] <= 77;
      opCodes[2267] <= 77;
      opCodes[2300] <= 77;
      opCodes[2308] <= 77;
      opCodes[2341] <= 77;
      opCodes[2393] <= 77;
      opCodes[2493] <= 77;
      opCodes[2504] <= 77;
      opCodes[2534] <= 77;
      opCodes[2545] <= 77;
      opCodes[2611] <= 77;
      opCodes[2646] <= 77;
      opCodes[2657] <= 77;
      opCodes[2687] <= 77;
      opCodes[2698] <= 77;
      opCodes[2728] <= 77;
      opCodes[2739] <= 77;
      opCodes[2787] <= 77;
      opCodes[2821] <= 77;
      opCodes[2937] <= 77;
      opCodes[2948] <= 77;
      opCodes[2975] <= 77;
      opCodes[2990] <= 77;
      opCodes[3027] <= 77;
      opCodes[152] <= 78;
      opCodes[226] <= 78;
      opCodes[822] <= 78;
      opCodes[896] <= 78;
      opCodes[1224] <= 78;
      opCodes[1298] <= 78;
      opCodes[153] <= 79;
      opCodes[227] <= 79;
      opCodes[230] <= 79;
      opCodes[823] <= 79;
      opCodes[897] <= 79;
      opCodes[900] <= 79;
      opCodes[1225] <= 79;
      opCodes[1299] <= 79;
      opCodes[1302] <= 79;
      opCodes[154] <= 80;
      opCodes[228] <= 80;
      opCodes[156] <= 81;
      opCodes[164] <= 81;
      opCodes[247] <= 81;
      opCodes[259] <= 81;
      opCodes[826] <= 81;
      opCodes[834] <= 81;
      opCodes[1228] <= 81;
      opCodes[1236] <= 81;
      opCodes[2870] <= 81;
      opCodes[2881] <= 81;
      opCodes[157] <= 82;
      opCodes[165] <= 82;
      opCodes[234] <= 82;
      opCodes[240] <= 82;
      opCodes[249] <= 82;
      opCodes[260] <= 82;
      opCodes[827] <= 82;
      opCodes[835] <= 82;
      opCodes[1229] <= 82;
      opCodes[1237] <= 82;
      opCodes[2871] <= 82;
      opCodes[2882] <= 82;
      opCodes[3061] <= 82;
      opCodes[158] <= 83;
      opCodes[160] <= 83;
      opCodes[241] <= 83;
      opCodes[243] <= 83;
      opCodes[828] <= 83;
      opCodes[830] <= 83;
      opCodes[1230] <= 83;
      opCodes[1232] <= 83;
      opCodes[1350] <= 83;
      opCodes[1352] <= 83;
      opCodes[1356] <= 83;
      opCodes[1358] <= 83;
      opCodes[2011] <= 83;
      opCodes[2013] <= 83;
      opCodes[2017] <= 83;
      opCodes[2019] <= 83;
      opCodes[2444] <= 83;
      opCodes[2446] <= 83;
      opCodes[2450] <= 83;
      opCodes[2452] <= 83;
      opCodes[159] <= 84;
      opCodes[242] <= 84;
      opCodes[829] <= 84;
      opCodes[1231] <= 84;
      opCodes[1351] <= 84;
      opCodes[1357] <= 84;
      opCodes[2012] <= 84;
      opCodes[2018] <= 84;
      opCodes[2445] <= 84;
      opCodes[2451] <= 84;
      opCodes[161] <= 85;
      opCodes[244] <= 85;
      opCodes[831] <= 85;
      opCodes[1233] <= 85;
      opCodes[1353] <= 85;
      opCodes[1359] <= 85;
      opCodes[2014] <= 85;
      opCodes[2020] <= 85;
      opCodes[2447] <= 85;
      opCodes[2453] <= 85;
      opCodes[162] <= 86;
      opCodes[245] <= 86;
      opCodes[832] <= 86;
      opCodes[1234] <= 86;
      opCodes[1366] <= 86;
      opCodes[1693] <= 86;
      opCodes[1840] <= 86;
      opCodes[2027] <= 86;
      opCodes[2302] <= 86;
      opCodes[2460] <= 86;
      opCodes[2700] <= 86;
      opCodes[163] <= 87;
      opCodes[246] <= 87;
      opCodes[258] <= 87;
      opCodes[833] <= 87;
      opCodes[1235] <= 87;
      opCodes[2880] <= 87;
      opCodes[166] <= 88;
      opCodes[176] <= 89;
      opCodes[189] <= 89;
      opCodes[178] <= 90;
      opCodes[184] <= 91;
      opCodes[190] <= 92;
      opCodes[198] <= 93;
      opCodes[868] <= 93;
      opCodes[1048] <= 93;
      opCodes[1270] <= 93;
      opCodes[3000] <= 93;
      opCodes[200] <= 94;
      opCodes[214] <= 94;
      opCodes[870] <= 94;
      opCodes[884] <= 94;
      opCodes[1050] <= 94;
      opCodes[1064] <= 94;
      opCodes[1272] <= 94;
      opCodes[1286] <= 94;
      opCodes[3002] <= 94;
      opCodes[3016] <= 94;
      opCodes[201] <= 95;
      opCodes[212] <= 95;
      opCodes[871] <= 95;
      opCodes[882] <= 95;
      opCodes[1051] <= 95;
      opCodes[1062] <= 95;
      opCodes[1273] <= 95;
      opCodes[1284] <= 95;
      opCodes[3003] <= 95;
      opCodes[3014] <= 95;
      opCodes[202] <= 96;
      opCodes[205] <= 96;
      opCodes[217] <= 96;
      opCodes[872] <= 96;
      opCodes[875] <= 96;
      opCodes[887] <= 96;
      opCodes[1052] <= 96;
      opCodes[1055] <= 96;
      opCodes[1067] <= 96;
      opCodes[1274] <= 96;
      opCodes[1277] <= 96;
      opCodes[1289] <= 96;
      opCodes[3004] <= 96;
      opCodes[3007] <= 96;
      opCodes[3019] <= 96;
      opCodes[203] <= 97;
      opCodes[215] <= 97;
      opCodes[873] <= 97;
      opCodes[885] <= 97;
      opCodes[1053] <= 97;
      opCodes[1065] <= 97;
      opCodes[1275] <= 97;
      opCodes[1287] <= 97;
      opCodes[3005] <= 97;
      opCodes[3017] <= 97;
      opCodes[206] <= 98;
      opCodes[876] <= 98;
      opCodes[1056] <= 98;
      opCodes[1278] <= 98;
      opCodes[3008] <= 98;
      opCodes[207] <= 99;
      opCodes[208] <= 100;
      opCodes[878] <= 100;
      opCodes[1058] <= 100;
      opCodes[1280] <= 100;
      opCodes[3010] <= 100;
      opCodes[209] <= 101;
      opCodes[879] <= 101;
      opCodes[1059] <= 101;
      opCodes[1281] <= 101;
      opCodes[3011] <= 101;
      opCodes[210] <= 102;
      opCodes[880] <= 102;
      opCodes[1060] <= 102;
      opCodes[1282] <= 102;
      opCodes[3012] <= 102;
      opCodes[211] <= 103;
      opCodes[881] <= 103;
      opCodes[1061] <= 103;
      opCodes[1283] <= 103;
      opCodes[3013] <= 103;
      opCodes[218] <= 104;
      opCodes[229] <= 105;
      opCodes[899] <= 105;
      opCodes[1301] <= 105;
      opCodes[231] <= 106;
      opCodes[901] <= 106;
      opCodes[232] <= 107;
      opCodes[902] <= 107;
      opCodes[233] <= 108;
      opCodes[239] <= 109;
      opCodes[248] <= 110;
      opCodes[250] <= 111;
      opCodes[252] <= 111;
      opCodes[255] <= 111;
      opCodes[1311] <= 111;
      opCodes[1314] <= 111;
      opCodes[1573] <= 111;
      opCodes[1575] <= 111;
      opCodes[1578] <= 111;
      opCodes[1582] <= 111;
      opCodes[1584] <= 111;
      opCodes[1587] <= 111;
      opCodes[1947] <= 111;
      opCodes[1949] <= 111;
      opCodes[1952] <= 111;
      opCodes[1969] <= 111;
      opCodes[1971] <= 111;
      opCodes[1974] <= 111;
      opCodes[2116] <= 111;
      opCodes[2118] <= 111;
      opCodes[2121] <= 111;
      opCodes[2125] <= 111;
      opCodes[2127] <= 111;
      opCodes[2130] <= 111;
      opCodes[2208] <= 111;
      opCodes[2210] <= 111;
      opCodes[2213] <= 111;
      opCodes[2549] <= 111;
      opCodes[2551] <= 111;
      opCodes[2554] <= 111;
      opCodes[2558] <= 111;
      opCodes[2560] <= 111;
      opCodes[2563] <= 111;
      opCodes[2872] <= 111;
      opCodes[2874] <= 111;
      opCodes[2877] <= 111;
      opCodes[251] <= 112;
      opCodes[1310] <= 112;
      opCodes[1574] <= 112;
      opCodes[1583] <= 112;
      opCodes[1948] <= 112;
      opCodes[1970] <= 112;
      opCodes[2117] <= 112;
      opCodes[2126] <= 112;
      opCodes[2209] <= 112;
      opCodes[2550] <= 112;
      opCodes[2559] <= 112;
      opCodes[2873] <= 112;
      opCodes[253] <= 113;
      opCodes[256] <= 113;
      opCodes[1312] <= 113;
      opCodes[1315] <= 113;
      opCodes[1576] <= 113;
      opCodes[1579] <= 113;
      opCodes[1585] <= 113;
      opCodes[1588] <= 113;
      opCodes[1950] <= 113;
      opCodes[1953] <= 113;
      opCodes[1972] <= 113;
      opCodes[1975] <= 113;
      opCodes[2119] <= 113;
      opCodes[2122] <= 113;
      opCodes[2128] <= 113;
      opCodes[2131] <= 113;
      opCodes[2211] <= 113;
      opCodes[2214] <= 113;
      opCodes[2552] <= 113;
      opCodes[2555] <= 113;
      opCodes[2561] <= 113;
      opCodes[2564] <= 113;
      opCodes[2875] <= 113;
      opCodes[2878] <= 113;
      opCodes[257] <= 114;
      opCodes[1598] <= 114;
      opCodes[2141] <= 114;
      opCodes[2574] <= 114;
      opCodes[2879] <= 114;
      opCodes[261] <= 115;
      opCodes[262] <= 116;
      opCodes[263] <= 117;
      opCodes[267] <= 118;
      opCodes[268] <= 119;
      opCodes[289] <= 119;
      opCodes[445] <= 119;
      opCodes[466] <= 119;
      opCodes[951] <= 119;
      opCodes[1550] <= 119;
      opCodes[1566] <= 119;
      opCodes[1916] <= 119;
      opCodes[1932] <= 119;
      opCodes[2354] <= 119;
      opCodes[2752] <= 119;
      opCodes[2890] <= 119;
      opCodes[269] <= 120;
      opCodes[270] <= 121;
      opCodes[286] <= 121;
      opCodes[337] <= 121;
      opCodes[393] <= 121;
      opCodes[419] <= 121;
      opCodes[271] <= 122;
      opCodes[273] <= 123;
      opCodes[274] <= 124;
      opCodes[295] <= 124;
      opCodes[451] <= 124;
      opCodes[472] <= 124;
      opCodes[957] <= 124;
      opCodes[1553] <= 124;
      opCodes[1569] <= 124;
      opCodes[1919] <= 124;
      opCodes[1935] <= 124;
      opCodes[2357] <= 124;
      opCodes[2755] <= 124;
      opCodes[2896] <= 124;
      opCodes[275] <= 125;
      opCodes[276] <= 126;
      opCodes[277] <= 127;
      opCodes[278] <= 128;
      opCodes[299] <= 128;
      opCodes[455] <= 128;
      opCodes[476] <= 128;
      opCodes[961] <= 128;
      opCodes[2900] <= 128;
      opCodes[279] <= 129;
      opCodes[300] <= 129;
      opCodes[456] <= 129;
      opCodes[477] <= 129;
      opCodes[962] <= 129;
      opCodes[2901] <= 129;
      opCodes[280] <= 130;
      opCodes[301] <= 130;
      opCodes[457] <= 130;
      opCodes[478] <= 130;
      opCodes[963] <= 130;
      opCodes[2902] <= 130;
      opCodes[281] <= 131;
      opCodes[302] <= 131;
      opCodes[458] <= 131;
      opCodes[479] <= 131;
      opCodes[964] <= 131;
      opCodes[2903] <= 131;
      opCodes[282] <= 132;
      opCodes[303] <= 132;
      opCodes[459] <= 132;
      opCodes[480] <= 132;
      opCodes[965] <= 132;
      opCodes[2904] <= 132;
      opCodes[283] <= 133;
      opCodes[304] <= 133;
      opCodes[460] <= 133;
      opCodes[481] <= 133;
      opCodes[966] <= 133;
      opCodes[2905] <= 133;
      opCodes[284] <= 134;
      opCodes[305] <= 134;
      opCodes[461] <= 134;
      opCodes[482] <= 134;
      opCodes[967] <= 134;
      opCodes[2906] <= 134;
      opCodes[285] <= 135;
      opCodes[306] <= 135;
      opCodes[462] <= 135;
      opCodes[483] <= 135;
      opCodes[968] <= 135;
      opCodes[2907] <= 135;
      opCodes[287] <= 136;
      opCodes[308] <= 136;
      opCodes[970] <= 136;
      opCodes[1536] <= 136;
      opCodes[288] <= 137;
      opCodes[309] <= 137;
      opCodes[971] <= 137;
      opCodes[1537] <= 137;
      opCodes[290] <= 138;
      opCodes[291] <= 139;
      opCodes[307] <= 139;
      opCodes[375] <= 139;
      opCodes[432] <= 139;
      opCodes[292] <= 140;
      opCodes[294] <= 141;
      opCodes[296] <= 142;
      opCodes[297] <= 143;
      opCodes[298] <= 144;
      opCodes[312] <= 145;
      opCodes[350] <= 145;
      opCodes[489] <= 145;
      opCodes[527] <= 145;
      opCodes[569] <= 145;
      opCodes[607] <= 145;
      opCodes[974] <= 145;
      opCodes[1376] <= 145;
      opCodes[1417] <= 145;
      opCodes[1458] <= 145;
      opCodes[1499] <= 145;
      opCodes[1615] <= 145;
      opCodes[1656] <= 145;
      opCodes[1697] <= 145;
      opCodes[1762] <= 145;
      opCodes[1803] <= 145;
      opCodes[1844] <= 145;
      opCodes[2469] <= 145;
      opCodes[2510] <= 145;
      opCodes[2622] <= 145;
      opCodes[2663] <= 145;
      opCodes[2704] <= 145;
      opCodes[2913] <= 145;
      opCodes[2951] <= 145;
      opCodes[318] <= 146;
      opCodes[356] <= 146;
      opCodes[495] <= 146;
      opCodes[533] <= 146;
      opCodes[575] <= 146;
      opCodes[613] <= 146;
      opCodes[980] <= 146;
      opCodes[1382] <= 146;
      opCodes[1423] <= 146;
      opCodes[1464] <= 146;
      opCodes[1505] <= 146;
      opCodes[1621] <= 146;
      opCodes[1662] <= 146;
      opCodes[1703] <= 146;
      opCodes[1768] <= 146;
      opCodes[1809] <= 146;
      opCodes[1850] <= 146;
      opCodes[2475] <= 146;
      opCodes[2516] <= 146;
      opCodes[2628] <= 146;
      opCodes[2669] <= 146;
      opCodes[2710] <= 146;
      opCodes[2919] <= 146;
      opCodes[2957] <= 146;
      opCodes[319] <= 147;
      opCodes[357] <= 147;
      opCodes[496] <= 147;
      opCodes[534] <= 147;
      opCodes[576] <= 147;
      opCodes[614] <= 147;
      opCodes[981] <= 147;
      opCodes[1383] <= 147;
      opCodes[1424] <= 147;
      opCodes[1465] <= 147;
      opCodes[1506] <= 147;
      opCodes[1622] <= 147;
      opCodes[1663] <= 147;
      opCodes[1704] <= 147;
      opCodes[1769] <= 147;
      opCodes[1810] <= 147;
      opCodes[1851] <= 147;
      opCodes[2476] <= 147;
      opCodes[2517] <= 147;
      opCodes[2629] <= 147;
      opCodes[2670] <= 147;
      opCodes[2711] <= 147;
      opCodes[2920] <= 147;
      opCodes[2958] <= 147;
      opCodes[320] <= 148;
      opCodes[358] <= 148;
      opCodes[497] <= 148;
      opCodes[535] <= 148;
      opCodes[577] <= 148;
      opCodes[615] <= 148;
      opCodes[982] <= 148;
      opCodes[1384] <= 148;
      opCodes[1425] <= 148;
      opCodes[1466] <= 148;
      opCodes[1507] <= 148;
      opCodes[1623] <= 148;
      opCodes[1664] <= 148;
      opCodes[1705] <= 148;
      opCodes[1770] <= 148;
      opCodes[1811] <= 148;
      opCodes[1852] <= 148;
      opCodes[2477] <= 148;
      opCodes[2518] <= 148;
      opCodes[2630] <= 148;
      opCodes[2671] <= 148;
      opCodes[2712] <= 148;
      opCodes[2921] <= 148;
      opCodes[2959] <= 148;
      opCodes[321] <= 149;
      opCodes[359] <= 149;
      opCodes[498] <= 149;
      opCodes[536] <= 149;
      opCodes[578] <= 149;
      opCodes[616] <= 149;
      opCodes[983] <= 149;
      opCodes[1385] <= 149;
      opCodes[1426] <= 149;
      opCodes[1467] <= 149;
      opCodes[1508] <= 149;
      opCodes[1624] <= 149;
      opCodes[1665] <= 149;
      opCodes[1706] <= 149;
      opCodes[1771] <= 149;
      opCodes[1812] <= 149;
      opCodes[1853] <= 149;
      opCodes[2478] <= 149;
      opCodes[2519] <= 149;
      opCodes[2631] <= 149;
      opCodes[2672] <= 149;
      opCodes[2713] <= 149;
      opCodes[2922] <= 149;
      opCodes[2960] <= 149;
      opCodes[322] <= 150;
      opCodes[323] <= 151;
      opCodes[361] <= 151;
      opCodes[500] <= 151;
      opCodes[538] <= 151;
      opCodes[580] <= 151;
      opCodes[618] <= 151;
      opCodes[985] <= 151;
      opCodes[1387] <= 151;
      opCodes[1428] <= 151;
      opCodes[1469] <= 151;
      opCodes[1510] <= 151;
      opCodes[1626] <= 151;
      opCodes[1667] <= 151;
      opCodes[1708] <= 151;
      opCodes[1773] <= 151;
      opCodes[1814] <= 151;
      opCodes[1855] <= 151;
      opCodes[2480] <= 151;
      opCodes[2521] <= 151;
      opCodes[2633] <= 151;
      opCodes[2674] <= 151;
      opCodes[2715] <= 151;
      opCodes[2924] <= 151;
      opCodes[2962] <= 151;
      opCodes[324] <= 152;
      opCodes[362] <= 152;
      opCodes[501] <= 152;
      opCodes[539] <= 152;
      opCodes[581] <= 152;
      opCodes[619] <= 152;
      opCodes[986] <= 152;
      opCodes[1388] <= 152;
      opCodes[1429] <= 152;
      opCodes[1470] <= 152;
      opCodes[1511] <= 152;
      opCodes[1627] <= 152;
      opCodes[1668] <= 152;
      opCodes[1709] <= 152;
      opCodes[1774] <= 152;
      opCodes[1815] <= 152;
      opCodes[1856] <= 152;
      opCodes[2481] <= 152;
      opCodes[2522] <= 152;
      opCodes[2634] <= 152;
      opCodes[2675] <= 152;
      opCodes[2716] <= 152;
      opCodes[2925] <= 152;
      opCodes[2963] <= 152;
      opCodes[325] <= 153;
      opCodes[363] <= 153;
      opCodes[502] <= 153;
      opCodes[540] <= 153;
      opCodes[582] <= 153;
      opCodes[620] <= 153;
      opCodes[987] <= 153;
      opCodes[1389] <= 153;
      opCodes[1430] <= 153;
      opCodes[1471] <= 153;
      opCodes[1512] <= 153;
      opCodes[1628] <= 153;
      opCodes[1669] <= 153;
      opCodes[1710] <= 153;
      opCodes[1775] <= 153;
      opCodes[1816] <= 153;
      opCodes[1857] <= 153;
      opCodes[2482] <= 153;
      opCodes[2523] <= 153;
      opCodes[2635] <= 153;
      opCodes[2676] <= 153;
      opCodes[2717] <= 153;
      opCodes[2926] <= 153;
      opCodes[2964] <= 153;
      opCodes[326] <= 154;
      opCodes[364] <= 154;
      opCodes[503] <= 154;
      opCodes[541] <= 154;
      opCodes[583] <= 154;
      opCodes[621] <= 154;
      opCodes[988] <= 154;
      opCodes[1390] <= 154;
      opCodes[1431] <= 154;
      opCodes[1472] <= 154;
      opCodes[1513] <= 154;
      opCodes[1629] <= 154;
      opCodes[1670] <= 154;
      opCodes[1711] <= 154;
      opCodes[1776] <= 154;
      opCodes[1817] <= 154;
      opCodes[1858] <= 154;
      opCodes[2483] <= 154;
      opCodes[2524] <= 154;
      opCodes[2636] <= 154;
      opCodes[2677] <= 154;
      opCodes[2718] <= 154;
      opCodes[2927] <= 154;
      opCodes[2965] <= 154;
      opCodes[327] <= 155;
      opCodes[365] <= 155;
      opCodes[504] <= 155;
      opCodes[542] <= 155;
      opCodes[584] <= 155;
      opCodes[622] <= 155;
      opCodes[989] <= 155;
      opCodes[1391] <= 155;
      opCodes[1432] <= 155;
      opCodes[1473] <= 155;
      opCodes[1514] <= 155;
      opCodes[1630] <= 155;
      opCodes[1671] <= 155;
      opCodes[1712] <= 155;
      opCodes[1777] <= 155;
      opCodes[1818] <= 155;
      opCodes[1859] <= 155;
      opCodes[2484] <= 155;
      opCodes[2525] <= 155;
      opCodes[2637] <= 155;
      opCodes[2678] <= 155;
      opCodes[2719] <= 155;
      opCodes[2928] <= 155;
      opCodes[2966] <= 155;
      opCodes[329] <= 156;
      opCodes[367] <= 156;
      opCodes[506] <= 156;
      opCodes[544] <= 156;
      opCodes[586] <= 156;
      opCodes[624] <= 156;
      opCodes[991] <= 156;
      opCodes[1393] <= 156;
      opCodes[1434] <= 156;
      opCodes[1475] <= 156;
      opCodes[1516] <= 156;
      opCodes[1632] <= 156;
      opCodes[1673] <= 156;
      opCodes[1714] <= 156;
      opCodes[1779] <= 156;
      opCodes[1820] <= 156;
      opCodes[1861] <= 156;
      opCodes[2486] <= 156;
      opCodes[2527] <= 156;
      opCodes[2639] <= 156;
      opCodes[2680] <= 156;
      opCodes[2721] <= 156;
      opCodes[2930] <= 156;
      opCodes[2968] <= 156;
      opCodes[330] <= 157;
      opCodes[368] <= 157;
      opCodes[507] <= 157;
      opCodes[545] <= 157;
      opCodes[587] <= 157;
      opCodes[625] <= 157;
      opCodes[992] <= 157;
      opCodes[1394] <= 157;
      opCodes[1435] <= 157;
      opCodes[1476] <= 157;
      opCodes[1517] <= 157;
      opCodes[1633] <= 157;
      opCodes[1674] <= 157;
      opCodes[1715] <= 157;
      opCodes[1780] <= 157;
      opCodes[1821] <= 157;
      opCodes[1862] <= 157;
      opCodes[2487] <= 157;
      opCodes[2528] <= 157;
      opCodes[2640] <= 157;
      opCodes[2681] <= 157;
      opCodes[2722] <= 157;
      opCodes[2931] <= 157;
      opCodes[2969] <= 157;
      opCodes[332] <= 158;
      opCodes[370] <= 158;
      opCodes[509] <= 158;
      opCodes[547] <= 158;
      opCodes[589] <= 158;
      opCodes[627] <= 158;
      opCodes[994] <= 158;
      opCodes[1396] <= 158;
      opCodes[1437] <= 158;
      opCodes[1478] <= 158;
      opCodes[1519] <= 158;
      opCodes[1635] <= 158;
      opCodes[1676] <= 158;
      opCodes[1717] <= 158;
      opCodes[1782] <= 158;
      opCodes[1823] <= 158;
      opCodes[1864] <= 158;
      opCodes[2489] <= 158;
      opCodes[2530] <= 158;
      opCodes[2642] <= 158;
      opCodes[2683] <= 158;
      opCodes[2724] <= 158;
      opCodes[2933] <= 158;
      opCodes[2971] <= 158;
      opCodes[333] <= 159;
      opCodes[360] <= 160;
      opCodes[371] <= 161;
      opCodes[392] <= 162;
      opCodes[405] <= 163;
      opCodes[406] <= 164;
      opCodes[407] <= 165;
      opCodes[409] <= 165;
      opCodes[412] <= 165;
      opCodes[408] <= 166;
      opCodes[410] <= 167;
      opCodes[417] <= 167;
      opCodes[411] <= 168;
      opCodes[1037] <= 168;
      opCodes[413] <= 169;
      opCodes[416] <= 170;
      opCodes[647] <= 170;
      opCodes[1370] <= 170;
      opCodes[1609] <= 170;
      opCodes[444] <= 171;
      opCodes[446] <= 172;
      opCodes[447] <= 173;
      opCodes[463] <= 173;
      opCodes[514] <= 173;
      opCodes[554] <= 173;
      opCodes[650] <= 173;
      opCodes[448] <= 174;
      opCodes[450] <= 175;
      opCodes[452] <= 176;
      opCodes[453] <= 177;
      opCodes[454] <= 178;
      opCodes[464] <= 179;
      opCodes[485] <= 179;
      opCodes[2909] <= 179;
      opCodes[465] <= 180;
      opCodes[486] <= 180;
      opCodes[2910] <= 180;
      opCodes[467] <= 181;
      opCodes[468] <= 182;
      opCodes[484] <= 182;
      opCodes[594] <= 182;
      opCodes[632] <= 182;
      opCodes[663] <= 182;
      opCodes[469] <= 183;
      opCodes[471] <= 184;
      opCodes[473] <= 185;
      opCodes[474] <= 186;
      opCodes[475] <= 187;
      opCodes[499] <= 188;
      opCodes[510] <= 189;
      opCodes[537] <= 190;
      opCodes[548] <= 191;
      opCodes[553] <= 192;
      opCodes[579] <= 193;
      opCodes[590] <= 194;
      opCodes[617] <= 195;
      opCodes[628] <= 196;
      opCodes[648] <= 197;
      opCodes[679] <= 198;
      opCodes[688] <= 199;
      opCodes[701] <= 199;
      opCodes[690] <= 200;
      opCodes[696] <= 201;
      opCodes[702] <= 202;
      opCodes[713] <= 203;
      opCodes[792] <= 203;
      opCodes[729] <= 204;
      opCodes[742] <= 204;
      opCodes[731] <= 205;
      opCodes[737] <= 206;
      opCodes[743] <= 207;
      opCodes[755] <= 208;
      opCodes[765] <= 209;
      opCodes[778] <= 209;
      opCodes[767] <= 210;
      opCodes[773] <= 211;
      opCodes[779] <= 212;
      opCodes[800] <= 213;
      opCodes[801] <= 214;
      opCodes[804] <= 215;
      opCodes[818] <= 216;
      opCodes[824] <= 217;
      opCodes[898] <= 217;
      opCodes[836] <= 218;
      opCodes[846] <= 219;
      opCodes[859] <= 219;
      opCodes[848] <= 220;
      opCodes[854] <= 221;
      opCodes[860] <= 222;
      opCodes[877] <= 223;
      opCodes[888] <= 224;
      opCodes[905] <= 225;
      opCodes[918] <= 226;
      opCodes[931] <= 226;
      opCodes[920] <= 227;
      opCodes[926] <= 228;
      opCodes[932] <= 229;
      opCodes[944] <= 230;
      opCodes[946] <= 231;
      opCodes[948] <= 232;
      opCodes[950] <= 233;
      opCodes[952] <= 234;
      opCodes[953] <= 235;
      opCodes[969] <= 235;
      opCodes[999] <= 235;
      opCodes[1019] <= 235;
      opCodes[1043] <= 235;
      opCodes[954] <= 236;
      opCodes[956] <= 237;
      opCodes[958] <= 238;
      opCodes[959] <= 239;
      opCodes[960] <= 240;
      opCodes[972] <= 241;
      opCodes[1010] <= 241;
      opCodes[984] <= 242;
      opCodes[995] <= 243;
      opCodes[1018] <= 244;
      opCodes[1031] <= 245;
      opCodes[1032] <= 246;
      opCodes[1033] <= 247;
      opCodes[1035] <= 247;
      opCodes[1038] <= 247;
      opCodes[1034] <= 248;
      opCodes[1036] <= 249;
      opCodes[1041] <= 249;
      opCodes[1039] <= 250;
      opCodes[1045] <= 251;
      opCodes[1057] <= 252;
      opCodes[1068] <= 253;
      opCodes[1081] <= 254;
      opCodes[1090] <= 255;
      opCodes[1103] <= 255;
      opCodes[1092] <= 256;
      opCodes[1098] <= 257;
      opCodes[1104] <= 258;
      opCodes[1115] <= 259;
      opCodes[1194] <= 259;
      opCodes[1131] <= 260;
      opCodes[1144] <= 260;
      opCodes[1133] <= 261;
      opCodes[1139] <= 262;
      opCodes[1145] <= 263;
      opCodes[1157] <= 264;
      opCodes[1167] <= 265;
      opCodes[1180] <= 265;
      opCodes[1169] <= 266;
      opCodes[1175] <= 267;
      opCodes[1181] <= 268;
      opCodes[1202] <= 269;
      opCodes[1203] <= 270;
      opCodes[1206] <= 271;
      opCodes[1220] <= 272;
      opCodes[1226] <= 273;
      opCodes[1300] <= 273;
      opCodes[1238] <= 274;
      opCodes[1248] <= 275;
      opCodes[1261] <= 275;
      opCodes[1250] <= 276;
      opCodes[1256] <= 277;
      opCodes[1262] <= 278;
      opCodes[1279] <= 279;
      opCodes[1290] <= 280;
      opCodes[1304] <= 281;
      opCodes[1308] <= 282;
      opCodes[1319] <= 282;
      opCodes[1367] <= 282;
      opCodes[1571] <= 282;
      opCodes[1599] <= 282;
      opCodes[1309] <= 283;
      opCodes[1316] <= 284;
      opCodes[1317] <= 285;
      opCodes[1318] <= 286;
      opCodes[1413] <= 286;
      opCodes[1495] <= 286;
      opCodes[1652] <= 286;
      opCodes[1799] <= 286;
      opCodes[2073] <= 286;
      opCodes[2261] <= 286;
      opCodes[2506] <= 286;
      opCodes[2659] <= 286;
      opCodes[1327] <= 287;
      opCodes[1338] <= 288;
      opCodes[1340] <= 289;
      opCodes[1346] <= 289;
      opCodes[2001] <= 289;
      opCodes[2007] <= 289;
      opCodes[2434] <= 289;
      opCodes[2440] <= 289;
      opCodes[1341] <= 290;
      opCodes[2002] <= 290;
      opCodes[2435] <= 290;
      opCodes[1347] <= 291;
      opCodes[1570] <= 291;
      opCodes[2008] <= 291;
      opCodes[2113] <= 291;
      opCodes[2441] <= 291;
      opCodes[2546] <= 291;
      opCodes[1348] <= 292;
      opCodes[1349] <= 293;
      opCodes[1374] <= 293;
      opCodes[1415] <= 293;
      opCodes[1538] <= 293;
      opCodes[1552] <= 293;
      opCodes[1572] <= 293;
      opCodes[1613] <= 293;
      opCodes[1654] <= 293;
      opCodes[1695] <= 293;
      opCodes[1733] <= 293;
      opCodes[1904] <= 293;
      opCodes[1918] <= 293;
      opCodes[1354] <= 294;
      opCodes[1580] <= 294;
      opCodes[1355] <= 295;
      opCodes[1456] <= 295;
      opCodes[1497] <= 295;
      opCodes[1554] <= 295;
      opCodes[1568] <= 295;
      opCodes[1581] <= 295;
      opCodes[1760] <= 295;
      opCodes[1801] <= 295;
      opCodes[1842] <= 295;
      opCodes[1880] <= 295;
      opCodes[1920] <= 295;
      opCodes[1934] <= 295;
      opCodes[1360] <= 296;
      opCodes[1589] <= 296;
      opCodes[1361] <= 297;
      opCodes[1371] <= 297;
      opCodes[1412] <= 297;
      opCodes[1590] <= 297;
      opCodes[1610] <= 297;
      opCodes[1651] <= 297;
      opCodes[1692] <= 297;
      opCodes[1362] <= 298;
      opCodes[1364] <= 298;
      opCodes[1591] <= 298;
      opCodes[1593] <= 298;
      opCodes[1596] <= 298;
      opCodes[1363] <= 299;
      opCodes[1592] <= 299;
      opCodes[1365] <= 300;
      opCodes[1594] <= 300;
      opCodes[1597] <= 300;
      opCodes[1372] <= 301;
      opCodes[1454] <= 301;
      opCodes[1611] <= 301;
      opCodes[1758] <= 301;
      opCodes[2032] <= 301;
      opCodes[2220] <= 301;
      opCodes[2465] <= 301;
      opCodes[2618] <= 301;
      opCodes[1373] <= 302;
      opCodes[1414] <= 302;
      opCodes[1386] <= 303;
      opCodes[1397] <= 304;
      opCodes[1427] <= 305;
      opCodes[1438] <= 306;
      opCodes[1453] <= 307;
      opCodes[1494] <= 307;
      opCodes[1757] <= 307;
      opCodes[1798] <= 307;
      opCodes[1839] <= 307;
      opCodes[1455] <= 308;
      opCodes[1496] <= 308;
      opCodes[1468] <= 309;
      opCodes[1479] <= 310;
      opCodes[1509] <= 311;
      opCodes[1520] <= 312;
      opCodes[1539] <= 313;
      opCodes[1905] <= 313;
      opCodes[1540] <= 314;
      opCodes[1906] <= 314;
      opCodes[1541] <= 315;
      opCodes[1907] <= 315;
      opCodes[1542] <= 316;
      opCodes[1558] <= 316;
      opCodes[1908] <= 316;
      opCodes[1924] <= 316;
      opCodes[2346] <= 316;
      opCodes[2744] <= 316;
      opCodes[1543] <= 317;
      opCodes[1559] <= 317;
      opCodes[1909] <= 317;
      opCodes[1925] <= 317;
      opCodes[2347] <= 317;
      opCodes[2745] <= 317;
      opCodes[1544] <= 318;
      opCodes[1560] <= 318;
      opCodes[1910] <= 318;
      opCodes[1926] <= 318;
      opCodes[2348] <= 318;
      opCodes[2746] <= 318;
      opCodes[1545] <= 319;
      opCodes[1561] <= 319;
      opCodes[1911] <= 319;
      opCodes[1927] <= 319;
      opCodes[2349] <= 319;
      opCodes[2747] <= 319;
      opCodes[1546] <= 320;
      opCodes[1562] <= 320;
      opCodes[1912] <= 320;
      opCodes[1928] <= 320;
      opCodes[2350] <= 320;
      opCodes[2748] <= 320;
      opCodes[1547] <= 321;
      opCodes[1563] <= 321;
      opCodes[1913] <= 321;
      opCodes[1929] <= 321;
      opCodes[2351] <= 321;
      opCodes[2749] <= 321;
      opCodes[1548] <= 322;
      opCodes[1564] <= 322;
      opCodes[1914] <= 322;
      opCodes[1930] <= 322;
      opCodes[2352] <= 322;
      opCodes[2750] <= 322;
      opCodes[1549] <= 323;
      opCodes[1565] <= 323;
      opCodes[1915] <= 323;
      opCodes[1931] <= 323;
      opCodes[2353] <= 323;
      opCodes[2751] <= 323;
      opCodes[1551] <= 324;
      opCodes[1917] <= 324;
      opCodes[1555] <= 325;
      opCodes[1921] <= 325;
      opCodes[1556] <= 326;
      opCodes[1922] <= 326;
      opCodes[1557] <= 327;
      opCodes[1923] <= 327;
      opCodes[1567] <= 328;
      opCodes[1933] <= 328;
      opCodes[1608] <= 329;
      opCodes[1612] <= 330;
      opCodes[1653] <= 330;
      opCodes[1694] <= 330;
      opCodes[1625] <= 331;
      opCodes[1636] <= 332;
      opCodes[1666] <= 333;
      opCodes[1677] <= 334;
      opCodes[1707] <= 335;
      opCodes[1718] <= 336;
      opCodes[1746] <= 337;
      opCodes[1759] <= 338;
      opCodes[1800] <= 338;
      opCodes[1841] <= 338;
      opCodes[1772] <= 339;
      opCodes[1783] <= 340;
      opCodes[1813] <= 341;
      opCodes[1824] <= 342;
      opCodes[1854] <= 343;
      opCodes[1865] <= 344;
      opCodes[1938] <= 345;
      opCodes[1939] <= 346;
      opCodes[1945] <= 347;
      opCodes[1954] <= 348;
      opCodes[1957] <= 348;
      opCodes[1955] <= 349;
      opCodes[1958] <= 350;
      opCodes[1959] <= 351;
      opCodes[1960] <= 352;
      opCodes[1962] <= 353;
      opCodes[1963] <= 354;
      opCodes[2397] <= 354;
      opCodes[2402] <= 354;
      opCodes[2823] <= 354;
      opCodes[1964] <= 355;
      opCodes[1965] <= 356;
      opCodes[1966] <= 357;
      opCodes[1981] <= 357;
      opCodes[1992] <= 357;
      opCodes[2145] <= 357;
      opCodes[2360] <= 357;
      opCodes[1967] <= 358;
      opCodes[1968] <= 359;
      opCodes[1979] <= 359;
      opCodes[2000] <= 359;
      opCodes[2143] <= 359;
      opCodes[2358] <= 359;
      opCodes[1976] <= 360;
      opCodes[1977] <= 361;
      opCodes[1978] <= 362;
      opCodes[2028] <= 362;
      opCodes[1991] <= 363;
      opCodes[1999] <= 364;
      opCodes[2009] <= 365;
      opCodes[2010] <= 366;
      opCodes[2034] <= 366;
      opCodes[2075] <= 366;
      opCodes[2115] <= 366;
      opCodes[2156] <= 366;
      opCodes[2196] <= 366;
      opCodes[2207] <= 366;
      opCodes[2222] <= 366;
      opCodes[2263] <= 366;
      opCodes[2304] <= 366;
      opCodes[2342] <= 366;
      opCodes[2356] <= 366;
      opCodes[2015] <= 367;
      opCodes[2123] <= 367;
      opCodes[2016] <= 368;
      opCodes[2045] <= 368;
      opCodes[2086] <= 368;
      opCodes[2124] <= 368;
      opCodes[2167] <= 368;
      opCodes[2233] <= 368;
      opCodes[2274] <= 368;
      opCodes[2315] <= 368;
      opCodes[2021] <= 369;
      opCodes[2132] <= 369;
      opCodes[2022] <= 370;
      opCodes[2133] <= 370;
      opCodes[2023] <= 371;
      opCodes[2025] <= 371;
      opCodes[2134] <= 371;
      opCodes[2137] <= 371;
      opCodes[2139] <= 371;
      opCodes[2024] <= 372;
      opCodes[2138] <= 372;
      opCodes[2026] <= 373;
      opCodes[2135] <= 373;
      opCodes[2140] <= 373;
      opCodes[2029] <= 374;
      opCodes[2030] <= 375;
      opCodes[2215] <= 375;
      opCodes[2218] <= 375;
      opCodes[2031] <= 376;
      opCodes[2072] <= 376;
      opCodes[2216] <= 376;
      opCodes[2219] <= 376;
      opCodes[2260] <= 376;
      opCodes[2301] <= 376;
      opCodes[2033] <= 377;
      opCodes[2074] <= 377;
      opCodes[2048] <= 378;
      opCodes[2062] <= 378;
      opCodes[2089] <= 378;
      opCodes[2103] <= 378;
      opCodes[2172] <= 378;
      opCodes[2186] <= 378;
      opCodes[2236] <= 378;
      opCodes[2250] <= 378;
      opCodes[2277] <= 378;
      opCodes[2291] <= 378;
      opCodes[2318] <= 378;
      opCodes[2332] <= 378;
      opCodes[2049] <= 379;
      opCodes[2051] <= 379;
      opCodes[2060] <= 379;
      opCodes[2090] <= 379;
      opCodes[2092] <= 379;
      opCodes[2101] <= 379;
      opCodes[2173] <= 379;
      opCodes[2175] <= 379;
      opCodes[2184] <= 379;
      opCodes[2237] <= 379;
      opCodes[2239] <= 379;
      opCodes[2248] <= 379;
      opCodes[2278] <= 379;
      opCodes[2280] <= 379;
      opCodes[2289] <= 379;
      opCodes[2319] <= 379;
      opCodes[2321] <= 379;
      opCodes[2330] <= 379;
      opCodes[2050] <= 380;
      opCodes[2052] <= 381;
      opCodes[2055] <= 381;
      opCodes[2093] <= 381;
      opCodes[2096] <= 381;
      opCodes[2176] <= 381;
      opCodes[2179] <= 381;
      opCodes[2240] <= 381;
      opCodes[2243] <= 381;
      opCodes[2281] <= 381;
      opCodes[2284] <= 381;
      opCodes[2322] <= 381;
      opCodes[2325] <= 381;
      opCodes[2053] <= 382;
      opCodes[2094] <= 382;
      opCodes[2177] <= 382;
      opCodes[2241] <= 382;
      opCodes[2282] <= 382;
      opCodes[2323] <= 382;
      opCodes[2056] <= 383;
      opCodes[2097] <= 383;
      opCodes[2180] <= 383;
      opCodes[2244] <= 383;
      opCodes[2285] <= 383;
      opCodes[2326] <= 383;
      opCodes[2057] <= 384;
      opCodes[2098] <= 384;
      opCodes[2181] <= 384;
      opCodes[2245] <= 384;
      opCodes[2286] <= 384;
      opCodes[2327] <= 384;
      opCodes[2058] <= 385;
      opCodes[2099] <= 385;
      opCodes[2182] <= 385;
      opCodes[2246] <= 385;
      opCodes[2287] <= 385;
      opCodes[2328] <= 385;
      opCodes[2059] <= 386;
      opCodes[2100] <= 386;
      opCodes[2183] <= 386;
      opCodes[2247] <= 386;
      opCodes[2288] <= 386;
      opCodes[2329] <= 386;
      opCodes[2063] <= 387;
      opCodes[2091] <= 388;
      opCodes[2104] <= 389;
      opCodes[2114] <= 390;
      opCodes[2142] <= 391;
      opCodes[2155] <= 392;
      opCodes[2169] <= 393;
      opCodes[2174] <= 394;
      opCodes[2187] <= 395;
      opCodes[2221] <= 396;
      opCodes[2262] <= 396;
      opCodes[2303] <= 396;
      opCodes[2238] <= 397;
      opCodes[2251] <= 398;
      opCodes[2279] <= 399;
      opCodes[2292] <= 400;
      opCodes[2320] <= 401;
      opCodes[2333] <= 402;
      opCodes[2343] <= 403;
      opCodes[2344] <= 404;
      opCodes[2345] <= 405;
      opCodes[2355] <= 406;
      opCodes[2366] <= 407;
      opCodes[2794] <= 407;
      opCodes[2368] <= 408;
      opCodes[2386] <= 408;
      opCodes[2796] <= 408;
      opCodes[2814] <= 408;
      opCodes[2369] <= 409;
      opCodes[2384] <= 409;
      opCodes[2797] <= 409;
      opCodes[2812] <= 409;
      opCodes[2370] <= 410;
      opCodes[2373] <= 410;
      opCodes[2389] <= 410;
      opCodes[2798] <= 410;
      opCodes[2801] <= 410;
      opCodes[2817] <= 410;
      opCodes[2371] <= 411;
      opCodes[2387] <= 411;
      opCodes[2799] <= 411;
      opCodes[2815] <= 411;
      opCodes[2378] <= 412;
      opCodes[2806] <= 412;
      opCodes[2379] <= 413;
      opCodes[2380] <= 414;
      opCodes[2808] <= 414;
      opCodes[2381] <= 415;
      opCodes[2809] <= 415;
      opCodes[2382] <= 416;
      opCodes[2810] <= 416;
      opCodes[2383] <= 417;
      opCodes[2811] <= 417;
      opCodes[2390] <= 418;
      opCodes[2394] <= 419;
      opCodes[2395] <= 420;
      opCodes[2396] <= 421;
      opCodes[2399] <= 422;
      opCodes[2825] <= 422;
      opCodes[2401] <= 423;
      opCodes[2403] <= 424;
      opCodes[2404] <= 425;
      opCodes[2405] <= 426;
      opCodes[2406] <= 427;
      opCodes[2409] <= 427;
      opCodes[2407] <= 428;
      opCodes[2410] <= 429;
      opCodes[2411] <= 430;
      opCodes[2412] <= 431;
      opCodes[2433] <= 431;
      opCodes[2589] <= 431;
      opCodes[2756] <= 431;
      opCodes[2414] <= 432;
      opCodes[2422] <= 432;
      opCodes[2591] <= 432;
      opCodes[2758] <= 432;
      opCodes[2769] <= 432;
      opCodes[2777] <= 432;
      opCodes[2788] <= 432;
      opCodes[2421] <= 433;
      opCodes[2432] <= 434;
      opCodes[2442] <= 435;
      opCodes[2443] <= 436;
      opCodes[2494] <= 436;
      opCodes[2535] <= 436;
      opCodes[2548] <= 436;
      opCodes[2576] <= 436;
      opCodes[2597] <= 436;
      opCodes[2647] <= 436;
      opCodes[2688] <= 436;
      opCodes[2729] <= 436;
      opCodes[2448] <= 437;
      opCodes[2556] <= 437;
      opCodes[2449] <= 438;
      opCodes[2467] <= 438;
      opCodes[2508] <= 438;
      opCodes[2557] <= 438;
      opCodes[2620] <= 438;
      opCodes[2661] <= 438;
      opCodes[2702] <= 438;
      opCodes[2740] <= 438;
      opCodes[2754] <= 438;
      opCodes[2454] <= 439;
      opCodes[2565] <= 439;
      opCodes[2455] <= 440;
      opCodes[2566] <= 440;
      opCodes[2601] <= 440;
      opCodes[2456] <= 441;
      opCodes[2458] <= 441;
      opCodes[2567] <= 441;
      opCodes[2570] <= 441;
      opCodes[2572] <= 441;
      opCodes[2457] <= 442;
      opCodes[2571] <= 442;
      opCodes[2459] <= 443;
      opCodes[2568] <= 443;
      opCodes[2573] <= 443;
      opCodes[2461] <= 444;
      opCodes[2575] <= 444;
      opCodes[2462] <= 445;
      opCodes[2463] <= 446;
      opCodes[2613] <= 446;
      opCodes[2616] <= 446;
      opCodes[2464] <= 447;
      opCodes[2505] <= 447;
      opCodes[2614] <= 447;
      opCodes[2617] <= 447;
      opCodes[2658] <= 447;
      opCodes[2699] <= 447;
      opCodes[2466] <= 448;
      opCodes[2507] <= 448;
      opCodes[2479] <= 449;
      opCodes[2490] <= 450;
      opCodes[2520] <= 451;
      opCodes[2531] <= 452;
      opCodes[2547] <= 453;
      opCodes[2588] <= 454;
      opCodes[2599] <= 455;
      opCodes[2608] <= 456;
      opCodes[2612] <= 457;
      opCodes[2619] <= 458;
      opCodes[2660] <= 458;
      opCodes[2701] <= 458;
      opCodes[2632] <= 459;
      opCodes[2643] <= 460;
      opCodes[2673] <= 461;
      opCodes[2684] <= 462;
      opCodes[2714] <= 463;
      opCodes[2725] <= 464;
      opCodes[2741] <= 465;
      opCodes[2742] <= 466;
      opCodes[2743] <= 467;
      opCodes[2753] <= 468;
      opCodes[2768] <= 469;
      opCodes[2775] <= 470;
      opCodes[2784] <= 471;
      opCodes[2807] <= 472;
      opCodes[2818] <= 473;
      opCodes[2822] <= 474;
      opCodes[2826] <= 475;
      opCodes[2829] <= 476;
      opCodes[2839] <= 477;
      opCodes[2852] <= 477;
      opCodes[2841] <= 478;
      opCodes[2847] <= 479;
      opCodes[2853] <= 480;
      opCodes[2860] <= 481;
      opCodes[2863] <= 481;
      opCodes[2862] <= 482;
      opCodes[2865] <= 483;
      opCodes[2866] <= 484;
      opCodes[2868] <= 485;
      opCodes[2883] <= 486;
      opCodes[2885] <= 487;
      opCodes[2887] <= 488;
      opCodes[2889] <= 489;
      opCodes[2891] <= 490;
      opCodes[2892] <= 491;
      opCodes[2908] <= 491;
      opCodes[2938] <= 491;
      opCodes[2978] <= 491;
      opCodes[2995] <= 491;
      opCodes[2893] <= 492;
      opCodes[2895] <= 493;
      opCodes[2897] <= 494;
      opCodes[2898] <= 495;
      opCodes[2899] <= 496;
      opCodes[2911] <= 497;
      opCodes[2949] <= 497;
      opCodes[2923] <= 498;
      opCodes[2934] <= 499;
      opCodes[2961] <= 500;
      opCodes[2972] <= 501;
      opCodes[2977] <= 502;
      opCodes[2991] <= 503;
      opCodes[2993] <= 504;
      opCodes[2997] <= 505;
      opCodes[3009] <= 506;
      opCodes[3020] <= 507;
      opCodes[3040] <= 508;
      opCodes[3053] <= 508;
      opCodes[3042] <= 509;
      opCodes[3048] <= 510;
      opCodes[3054] <= 511;
      opCodes[3062] <= 512;
      opCodes[3065] <= 513;
      opCodes[3068] <= 513;
      opCodes[3067] <= 514;
      opCodes[3070] <= 515;
      opCodes[3071] <= 516;

      memory[285] <= 4; /* put key*/
      memory[107] <= 4; /* put data */
    end
    else begin                                                                  // Run
      //$display("%4d %4d %4d s=%4d f=%4d d=%4d", steps, step, intermediateValue, stop, found, data);
      case(opCodes[step])
           0 : begin intermediateValue <= memory[285]/*put_Key*/; /* get 1 */ step <= step + 1; end
           1 : begin memory[111]/*findAndInsert_Key*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
           2 : begin intermediateValue <= memory[284]/*put_Data*/; /* get 1 */ step <= step + 1; end
           3 : begin memory[110]/*findAndInsert_Data*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
           4 : begin intermediateValue <= memory[111]/*findAndInsert_Key*/; /* get 1 */ step <= step + 1; end
           5 : begin memory[113]/*find_Key*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
           6 : begin intermediateValue <= memory[145+memory[287]/*root*/]/*isLeaf[root]*/; /* get 2 */ step <= step + 1; end
           7 : begin memory[288]/*rootIsLeaf*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
           8 : begin intermediateValue <= memory[288]/*rootIsLeaf*/; /* get 1 */ step <= step + 1; end
           9 : begin if (intermediateValue == 0) step <=   44; else step = step + 1;/* endIfEq*/    end
          10 : begin memory[348]/*stuck*/ <= 0; /* set 1 */ step <= step + 1; end
          11 : begin intermediateValue <= memory[113]/*find_Key*/; /* get 1 */ step <= step + 1; end
          12 : begin memory[294]/*s_key*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          13 : begin memory[292]/*s_found*/ <= 0; /* set 1 */ step <= step + 1; end
          14 : begin memory[293]/*s_index*/ <= 0; /* set 1 */ step <= step + 1; end
          15 : begin intermediateValue <= memory[5+memory[348]/*stuck*/]/*current_size[stuck]*/; /* get 2 */ step <= step + 1; end
          16 : begin memory[344]/*stuckSearch_N*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          17 : begin intermediateValue <= memory[293]/*s_index*/ < memory[344]/*stuckSearch_N*/ ? -1 : memory[293]/*s_index*/ == memory[344]/*stuckSearch_N*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
          18 : begin if (intermediateValue >= 0) step <=   33; else step = step + 1;/* endIfGe*/    end
          19 : begin intermediateValue <= memory[294]/*s_key*/ < memory[166+memory[348]/*stuck*/*4+memory[293]/*s_index*/]/*keys[s_index,stuck]*/ ? -1 : memory[294]/*s_key*/ == memory[166+memory[348]/*stuck*/*4+memory[293]/*s_index*/]/*keys[s_index,stuck]*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
          20 : begin if (intermediateValue != 0) step <=   27; else step = step + 1;/* endIfNe*/    end
          21 : begin memory[292]/*s_found*/ <= 1; /* set 1 */ step <= step + 1; end
          22 : begin intermediateValue <= memory[166+memory[348]/*stuck*/*4+memory[293]/*s_index*/]/*keys[s_index,stuck]*/; /* get 3 */ step <= step + 1; end
          23 : begin intermediateValue <= memory[25+memory[348]/*stuck*/*4+memory[293]/*s_index*/]/*data[s_index,stuck]*/; /* get 3 */ step <= step + 1; end
          24 : begin memory[289]/*s_data*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          25 : begin step <=   33; /* end */ end
          26 : begin intermediateValue <= memory[293]/*s_index*/; /* get 1 */ step <= step + 1; end
          27 : begin intermediateValue <= 1 + intermediateValue;  /* add 1 */ step <= step + 1; end
          28 : begin memory[293]/*s_index*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          29 : begin step <= 17; /* start */ end
          30 : begin intermediateValue <= memory[287]/*root*/; /* get 1 */ step <= step + 1; end
          31 : begin memory[118]/*f_leaf*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          32 : begin intermediateValue <= memory[292]/*s_found*/; /* get 1 */ step <= step + 1; end
          33 : begin memory[108]/*f_found*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          34 : begin memory[112]/*f_index*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          35 : begin intermediateValue <= memory[294]/*s_key*/; /* get 1 */ step <= step + 1; end
          36 : begin memory[117]/*f_key*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          37 : begin intermediateValue <= memory[289]/*s_data*/; /* get 1 */ step <= step + 1; end
          38 : begin memory[107]/*f_data*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          39 : begin step <=   133; /* end */ end
          40 : begin memory[283]/*parent*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          41 : begin memory[114] <= 0; /* clear 1 */ step <= step + 1; end
          42 : begin intermediateValue <= memory[283]/*parent*/; /* get 1 */ step <= step + 1; end
          43 : begin memory[348]/*stuck*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          44 : begin intermediateValue <= memory[344]/*stuckSearch_N*/; /* get 1 */ step <= step + 1; end
          45 : begin intermediateValue <= -1 + intermediateValue;  /* add 1 */ step <= step + 1; end
          46 : begin if (intermediateValue >= 0) step <=   74; else step = step + 1;/* endIfGe*/    end
          47 : begin if (intermediateValue >  0) step <=   68; else step = step + 1;/* endIfGt*/    end
          48 : begin step <=   74; /* end */ end
          49 : begin step <= 58; /* start */ end
          50 : begin memory[4]/*child*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          51 : begin intermediateValue <= memory[4]/*child*/; /* get 1 */ step <= step + 1; end
          52 : begin memory[142]/*isALeaf*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          53 : begin intermediateValue <= memory[145+memory[142]/*isALeaf*/]/*isLeaf[isALeaf]*/; /* get 2 */ step <= step + 1; end
          54 : begin intermediateValue <= memory[142]/*isALeaf*/; /* get 1 */ step <= step + 1; end
          55 : begin if (intermediateValue == 0) step <=   123; else step = step + 1;/* endIfEq*/    end
          56 : begin if (intermediateValue >= 0) step <=   110; else step = step + 1;/* endIfGe*/    end
          57 : begin if (intermediateValue != 0) step <=   104; else step = step + 1;/* endIfNe*/    end
          58 : begin step <=   110; /* end */ end
          59 : begin step <= 94; /* start */ end
          60 : begin memory[115]/*find_result_leaf*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          61 : begin intermediateValue <= memory[115]/*find_result_leaf*/; /* get 1 */ step <= step + 1; end
          62 : begin intermediateValue <= memory[114]/*find_loop*/; /* get 1 */ step <= step + 1; end
          63 : begin memory[114]/*find_loop*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          64 : begin intermediateValue <= 9 <  intermediateValue ? -1 : 9 == intermediateValue ?  0 : +1; /* compare 1 */ step <= step + 1; end
          65 : begin if (intermediateValue >= 0) step <=   132; else step = step + 1;/* endIfGe*/    end
          66 : begin step <= 47; /* start */ end
          67 : begin stopped <= 1; end
          68 : begin intermediateValue <= memory[108]/*f_found*/; /* get 1 */ step <= step + 1; end
          69 : begin if (intermediateValue == 0) step <=   155; else step = step + 1;/* endIfEq*/    end
          70 : begin intermediateValue <= memory[118]/*f_leaf*/; /* get 1 */ step <= step + 1; end
          71 : begin intermediateValue <= memory[110]/*findAndInsert_Data*/; /* get 1 */ step <= step + 1; end
          72 : begin intermediateValue <= memory[112]/*f_index*/; /* get 1 */ step <= step + 1; end
          73 : begin memory[166+memory[348]/*stuck*/*4+memory[293]/*s_index*/]/*keys[s_index,stuck]*/ <= intermediateValue; /* set 3 */ step <= step + 1; end
          74 : begin memory[25+memory[348]/*stuck*/*4+memory[293]/*s_index*/]/*data[s_index,stuck]*/ <= intermediateValue; /* set 3 */ step <= step + 1; end
          75 : begin intermediateValue <= memory[293]/*s_index*/ < memory[5+memory[348]/*stuck*/]/*current_size[stuck]*/ ? -1 : memory[293]/*s_index*/ == memory[5+memory[348]/*stuck*/]/*current_size[stuck]*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
          76 : begin if (intermediateValue <  0) step <=   152; else step = step + 1;/* endIfLt*/    end
          77 : begin memory[5+memory[348]/*stuck*/]/*current_size[stuck]*/ <= intermediateValue; /* set 2 */ step <= step + 1; end
          78 : begin memory[140]/*f_success*/ <= 1; /* set 1 */ step <= step + 1; end
          79 : begin memory[116]/*f_inserted*/ <= 0; /* set 1 */ step <= step + 1; end
          80 : begin step <=   231; /* end */ end
          81 : begin memory[144]/*isFull*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          82 : begin intermediateValue <= memory[144]/*isFull*/; /* get 1 */ step <= step + 1; end
          83 : begin memory[246]/*leafSize*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          84 : begin intermediateValue <= memory[5+memory[246]/*leafSize*/]/*current_size[leafSize]*/; /* get 2 */ step <= step + 1; end
          85 : begin intermediateValue <= memory[246]/*leafSize*/; /* get 1 */ step <= step + 1; end
          86 : begin intermediateValue <= 2 <  intermediateValue ? -1 : 2 == intermediateValue ?  0 : +1; /* compare 1 */ step <= step + 1; end
          87 : begin intermediateValue <= intermediateValue >= 0 ? 1 : 0; /* ge */ step <= step + 1; end
          88 : begin if (intermediateValue >  0) step <=   229; else step = step + 1;/* endIfGt*/    end
          89 : begin if (intermediateValue >= 0) step <=   191; else step = step + 1;/* endIfGe*/    end
          90 : begin if (intermediateValue >  0) step <=   185; else step = step + 1;/* endIfGt*/    end
          91 : begin step <=   191; /* end */ end
          92 : begin step <= 175; /* start */ end
          93 : begin memory[340]/*stuckInsertElementAt_L*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          94 : begin memory[339]/*stuckInsertElementAt_i*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          95 : begin intermediateValue <= memory[339]/*stuckInsertElementAt_i*/; /* get 1 */ step <= step + 1; end
          96 : begin memory[338]/*stuckInsertElementAt_I*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          97 : begin intermediateValue <= memory[338]/*stuckInsertElementAt_I*/; /* get 1 */ step <= step + 1; end
          98 : begin intermediateValue <= memory[339]/*stuckInsertElementAt_i*/ < memory[340]/*stuckInsertElementAt_L*/ ? -1 : memory[339]/*stuckInsertElementAt_i*/ == memory[340]/*stuckInsertElementAt_L*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
          99 : begin if (intermediateValue == 0) step <=   219; else step = step + 1;/* endIfEq*/    end
         100 : begin intermediateValue <= memory[166+memory[348]/*stuck*/*4+memory[338]/*stuckInsertElementAt_I*/]/*keys[stuckInsertElementAt_I,stuck]*/; /* get 3 */ step <= step + 1; end
         101 : begin memory[166+memory[348]/*stuck*/*4+memory[339]/*stuckInsertElementAt_i*/]/*keys[stuckInsertElementAt_i,stuck]*/ <= intermediateValue; /* set 3 */ step <= step + 1; end
         102 : begin intermediateValue <= memory[25+memory[348]/*stuck*/*4+memory[338]/*stuckInsertElementAt_I*/]/*data[stuckInsertElementAt_I,stuck]*/; /* get 3 */ step <= step + 1; end
         103 : begin memory[25+memory[348]/*stuck*/*4+memory[339]/*stuckInsertElementAt_i*/]/*data[stuckInsertElementAt_i,stuck]*/ <= intermediateValue; /* set 3 */ step <= step + 1; end
         104 : begin step <= 206; /* start */ end
         105 : begin memory[140]/*f_success*/ <= 0; /* set 1 */ step <= step + 1; end
         106 : begin intermediateValue <= memory[140]/*f_success*/; /* get 1 */ step <= step + 1; end
         107 : begin if (intermediateValue >  0) step <=   3073; else step = step + 1;/* endIfGt*/    end
         108 : begin memory[144] <= 0; /* clear 1 */ step <= step + 1; end
         109 : begin if (intermediateValue == 0) step <=   248; else step = step + 1;/* endIfEq*/    end
         110 : begin if (intermediateValue >  0) step <=   260; else step = step + 1;/* endIfGt*/    end
         111 : begin memory[3]/*branchSize*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         112 : begin intermediateValue <= memory[5+memory[3]/*branchSize*/]/*current_size[branchSize]*/; /* get 2 */ step <= step + 1; end
         113 : begin intermediateValue <= memory[3]/*branchSize*/; /* get 1 */ step <= step + 1; end
         114 : begin intermediateValue <= 3 <  intermediateValue ? -1 : 3 == intermediateValue ?  0 : +1; /* compare 1 */ step <= step + 1; end
         115 : begin memory[143]/*isFullRoot*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         116 : begin intermediateValue <= memory[143]/*isFullRoot*/; /* get 1 */ step <= step + 1; end
         117 : begin if (intermediateValue == 0) step <=   903; else step = step + 1;/* endIfEq*/    end
         118 : begin if (intermediateValue == 0) step <=   443; else step = step + 1;/* endIfEq*/    end
         119 : begin intermediateValue <= memory[119]/*freeChainHead*/; /* get 1 */ step <= step + 1; end
         120 : begin memory[314]/*splitLeafRoot_l*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         121 : begin intermediateValue <= memory[314]/*splitLeafRoot_l*/; /* get 1 */ step <= step + 1; end
         122 : begin if (intermediateValue >  0) step <=   273; else step = step + 1;/* endIfGt*/    end
         123 : begin intermediateValue <= memory[120+memory[314]/*splitLeafRoot_l*/]/*free[splitLeafRoot_l]*/; /* get 2 */ step <= step + 1; end
         124 : begin memory[119]/*freeChainHead*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         125 : begin memory[120+memory[314]/*splitLeafRoot_l*/]/*free[splitLeafRoot_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         126 : begin memory[145+memory[314]/*splitLeafRoot_l*/]/*isLeaf[splitLeafRoot_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         127 : begin memory[5+memory[314]/*splitLeafRoot_l*/]/*current_size[splitLeafRoot_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         128 : begin memory[166] <= 0; /* clear 2 */ step <= step + 1; end
         129 : begin memory[167] <= 0; /* clear 2 */ step <= step + 1; end
         130 : begin memory[168] <= 0; /* clear 2 */ step <= step + 1; end
         131 : begin memory[169] <= 0; /* clear 2 */ step <= step + 1; end
         132 : begin memory[25] <= 0; /* clear 2 */ step <= step + 1; end
         133 : begin memory[26] <= 0; /* clear 2 */ step <= step + 1; end
         134 : begin memory[27] <= 0; /* clear 2 */ step <= step + 1; end
         135 : begin memory[28] <= 0; /* clear 2 */ step <= step + 1; end
         136 : begin memory[291]/*setLeaf*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         137 : begin memory[145+memory[291]/*setLeaf*/]/*isLeaf[setLeaf]*/ <= 1; /* set 2 */ step <= step + 1; end
         138 : begin memory[315]/*splitLeafRoot_r*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         139 : begin intermediateValue <= memory[315]/*splitLeafRoot_r*/; /* get 1 */ step <= step + 1; end
         140 : begin if (intermediateValue >  0) step <=   294; else step = step + 1;/* endIfGt*/    end
         141 : begin intermediateValue <= memory[120+memory[315]/*splitLeafRoot_r*/]/*free[splitLeafRoot_r]*/; /* get 2 */ step <= step + 1; end
         142 : begin memory[120+memory[315]/*splitLeafRoot_r*/]/*free[splitLeafRoot_r]*/ <= 0; /* set 2 */ step <= step + 1; end
         143 : begin memory[145+memory[315]/*splitLeafRoot_r*/]/*isLeaf[splitLeafRoot_r]*/ <= 0; /* set 2 */ step <= step + 1; end
         144 : begin memory[5+memory[315]/*splitLeafRoot_r*/]/*current_size[splitLeafRoot_r]*/ <= 0; /* set 2 */ step <= step + 1; end
         145 : begin memory[293] <= 0; /* clear 1 */ step <= step + 1; end
         146 : begin memory[347]/*stuckShift_N*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         147 : begin memory[345]/*stuckShift_i*/ <= 0; /* set 1 */ step <= step + 1; end
         148 : begin memory[346]/*stuckShift_I*/ <= 1; /* set 1 */ step <= step + 1; end
         149 : begin intermediateValue <= memory[346]/*stuckShift_I*/ < memory[347]/*stuckShift_N*/ ? -1 : memory[346]/*stuckShift_I*/ == memory[347]/*stuckShift_N*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
         150 : begin if (intermediateValue >= 0) step <=   334; else step = step + 1;/* endIfGe*/    end
         151 : begin intermediateValue <= memory[166+memory[348]/*stuck*/*4+memory[346]/*stuckShift_I*/]/*keys[stuckShift_I,stuck]*/; /* get 3 */ step <= step + 1; end
         152 : begin memory[166+memory[348]/*stuck*/*4+memory[345]/*stuckShift_i*/]/*keys[stuckShift_i,stuck]*/ <= intermediateValue; /* set 3 */ step <= step + 1; end
         153 : begin intermediateValue <= memory[25+memory[348]/*stuck*/*4+memory[346]/*stuckShift_I*/]/*data[stuckShift_I,stuck]*/; /* get 3 */ step <= step + 1; end
         154 : begin memory[25+memory[348]/*stuck*/*4+memory[345]/*stuckShift_i*/]/*data[stuckShift_i,stuck]*/ <= intermediateValue; /* set 3 */ step <= step + 1; end
         155 : begin intermediateValue <= memory[345]/*stuckShift_i*/; /* get 1 */ step <= step + 1; end
         156 : begin memory[345]/*stuckShift_i*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         157 : begin intermediateValue <= memory[346]/*stuckShift_I*/; /* get 1 */ step <= step + 1; end
         158 : begin memory[346]/*stuckShift_I*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         159 : begin step <= 321; /* start */ end
         160 : begin if (intermediateValue >= 0) step <=   372; else step = step + 1;/* endIfGe*/    end
         161 : begin step <= 359; /* start */ end
         162 : begin memory[310]/*splitLeafRoot_first*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         163 : begin memory[313]/*splitLeafRoot_last*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         164 : begin intermediateValue <= memory[313]/*splitLeafRoot_last*/; /* get 1 */ step <= step + 1; end
         165 : begin memory[312]/*splitLeafRoot_kv*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         166 : begin intermediateValue <= memory[310]/*splitLeafRoot_first*/ + memory[312]/*splitLeafRoot_kv*/; /* add2 */ step <= step + 1; end
         167 : begin intermediateValue <= memory[312]/*splitLeafRoot_kv*/; /* get 1 */ step <= step + 1; end
         168 : begin intermediateValue <= intermediateValue >> 1; /* shift right */ step <= step + 1; end
         169 : begin memory[145+memory[287]/*root*/]/*isLeaf[root]*/ <= 0; /* set 2 */ step <= step + 1; end
         170 : begin memory[5+memory[348]/*stuck*/]/*current_size[stuck]*/ <= 0; /* set 2 */ step <= step + 1; end
         171 : begin if (intermediateValue >  0) step <=   674; else step = step + 1;/* endIfGt*/    end
         172 : begin memory[300]/*splitBranchRoot_l*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         173 : begin intermediateValue <= memory[300]/*splitBranchRoot_l*/; /* get 1 */ step <= step + 1; end
         174 : begin if (intermediateValue >  0) step <=   450; else step = step + 1;/* endIfGt*/    end
         175 : begin intermediateValue <= memory[120+memory[300]/*splitBranchRoot_l*/]/*free[splitBranchRoot_l]*/; /* get 2 */ step <= step + 1; end
         176 : begin memory[120+memory[300]/*splitBranchRoot_l*/]/*free[splitBranchRoot_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         177 : begin memory[145+memory[300]/*splitBranchRoot_l*/]/*isLeaf[splitBranchRoot_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         178 : begin memory[5+memory[300]/*splitBranchRoot_l*/]/*current_size[splitBranchRoot_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         179 : begin memory[290]/*setBranch*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         180 : begin memory[145+memory[290]/*setBranch*/]/*isLeaf[setBranch]*/ <= 0; /* set 2 */ step <= step + 1; end
         181 : begin memory[302]/*splitBranchRoot_r*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         182 : begin intermediateValue <= memory[302]/*splitBranchRoot_r*/; /* get 1 */ step <= step + 1; end
         183 : begin if (intermediateValue >  0) step <=   471; else step = step + 1;/* endIfGt*/    end
         184 : begin intermediateValue <= memory[120+memory[302]/*splitBranchRoot_r*/]/*free[splitBranchRoot_r]*/; /* get 2 */ step <= step + 1; end
         185 : begin memory[120+memory[302]/*splitBranchRoot_r*/]/*free[splitBranchRoot_r]*/ <= 0; /* set 2 */ step <= step + 1; end
         186 : begin memory[145+memory[302]/*splitBranchRoot_r*/]/*isLeaf[splitBranchRoot_r]*/ <= 0; /* set 2 */ step <= step + 1; end
         187 : begin memory[5+memory[302]/*splitBranchRoot_r*/]/*current_size[splitBranchRoot_r]*/ <= 0; /* set 2 */ step <= step + 1; end
         188 : begin if (intermediateValue >= 0) step <=   511; else step = step + 1;/* endIfGe*/    end
         189 : begin step <= 498; /* start */ end
         190 : begin if (intermediateValue >= 0) step <=   549; else step = step + 1;/* endIfGe*/    end
         191 : begin step <= 536; /* start */ end
         192 : begin memory[301]/*splitBranchRoot_plk*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         193 : begin if (intermediateValue >= 0) step <=   591; else step = step + 1;/* endIfGe*/    end
         194 : begin step <= 578; /* start */ end
         195 : begin if (intermediateValue >= 0) step <=   629; else step = step + 1;/* endIfGe*/    end
         196 : begin step <= 616; /* start */ end
         197 : begin intermediateValue <= memory[301]/*splitBranchRoot_plk*/; /* get 1 */ step <= step + 1; end
         198 : begin if (intermediateValue == 0) step <=   714; else step = step + 1;/* endIfEq*/    end
         199 : begin if (intermediateValue >= 0) step <=   703; else step = step + 1;/* endIfGe*/    end
         200 : begin if (intermediateValue != 0) step <=   697; else step = step + 1;/* endIfNe*/    end
         201 : begin step <=   703; /* end */ end
         202 : begin step <= 687; /* start */ end
         203 : begin step <=   803; /* end */ end
         204 : begin if (intermediateValue >= 0) step <=   744; else step = step + 1;/* endIfGe*/    end
         205 : begin if (intermediateValue >  0) step <=   738; else step = step + 1;/* endIfGt*/    end
         206 : begin step <=   744; /* end */ end
         207 : begin step <= 728; /* start */ end
         208 : begin if (intermediateValue == 0) step <=   793; else step = step + 1;/* endIfEq*/    end
         209 : begin if (intermediateValue >= 0) step <=   780; else step = step + 1;/* endIfGe*/    end
         210 : begin if (intermediateValue != 0) step <=   774; else step = step + 1;/* endIfNe*/    end
         211 : begin step <=   780; /* end */ end
         212 : begin step <= 764; /* start */ end
         213 : begin if (intermediateValue >= 0) step <=   802; else step = step + 1;/* endIfGe*/    end
         214 : begin step <= 717; /* start */ end
         215 : begin if (intermediateValue == 0) step <=   825; else step = step + 1;/* endIfEq*/    end
         216 : begin if (intermediateValue <  0) step <=   822; else step = step + 1;/* endIfLt*/    end
         217 : begin step <=   901; /* end */ end
         218 : begin if (intermediateValue >  0) step <=   899; else step = step + 1;/* endIfGt*/    end
         219 : begin if (intermediateValue >= 0) step <=   861; else step = step + 1;/* endIfGe*/    end
         220 : begin if (intermediateValue >  0) step <=   855; else step = step + 1;/* endIfGt*/    end
         221 : begin step <=   861; /* end */ end
         222 : begin step <= 845; /* start */ end
         223 : begin if (intermediateValue == 0) step <=   889; else step = step + 1;/* endIfEq*/    end
         224 : begin step <= 876; /* start */ end
         225 : begin memory[286] <= 0; /* clear 1 */ step <= step + 1; end
         226 : begin if (intermediateValue >= 0) step <=   933; else step = step + 1;/* endIfGe*/    end
         227 : begin if (intermediateValue >  0) step <=   927; else step = step + 1;/* endIfGt*/    end
         228 : begin step <=   933; /* end */ end
         229 : begin step <= 917; /* start */ end
         230 : begin if (intermediateValue == 0) step <=   2869; else step = step + 1;/* endIfEq*/    end
         231 : begin memory[308]/*splitLeaf_node*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         232 : begin memory[309]/*splitLeaf_parent*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         233 : begin memory[305]/*splitLeaf_index*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         234 : begin memory[307]/*splitLeaf_l*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         235 : begin intermediateValue <= memory[307]/*splitLeaf_l*/; /* get 1 */ step <= step + 1; end
         236 : begin if (intermediateValue >  0) step <=   956; else step = step + 1;/* endIfGt*/    end
         237 : begin intermediateValue <= memory[120+memory[307]/*splitLeaf_l*/]/*free[splitLeaf_l]*/; /* get 2 */ step <= step + 1; end
         238 : begin memory[120+memory[307]/*splitLeaf_l*/]/*free[splitLeaf_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         239 : begin memory[145+memory[307]/*splitLeaf_l*/]/*isLeaf[splitLeaf_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         240 : begin memory[5+memory[307]/*splitLeaf_l*/]/*current_size[splitLeaf_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         241 : begin intermediateValue <= memory[308]/*splitLeaf_node*/; /* get 1 */ step <= step + 1; end
         242 : begin if (intermediateValue >= 0) step <=   996; else step = step + 1;/* endIfGe*/    end
         243 : begin step <= 983; /* start */ end
         244 : begin memory[303]/*splitLeaf_F*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         245 : begin memory[306]/*splitLeaf_L*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         246 : begin intermediateValue <= memory[303]/*splitLeaf_F*/; /* get 1 */ step <= step + 1; end
         247 : begin memory[304]/*splitLeaf_fl*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         248 : begin intermediateValue <= memory[306]/*splitLeaf_L*/ + memory[304]/*splitLeaf_fl*/; /* add2 */ step <= step + 1; end
         249 : begin intermediateValue <= memory[304]/*splitLeaf_fl*/; /* get 1 */ step <= step + 1; end
         250 : begin intermediateValue <= memory[309]/*splitLeaf_parent*/; /* get 1 */ step <= step + 1; end
         251 : begin intermediateValue <= memory[305]/*splitLeaf_index*/; /* get 1 */ step <= step + 1; end
         252 : begin if (intermediateValue == 0) step <=   1069; else step = step + 1;/* endIfEq*/    end
         253 : begin step <= 1056; /* start */ end
         254 : begin if (intermediateValue == 0) step <=   1116; else step = step + 1;/* endIfEq*/    end
         255 : begin if (intermediateValue >= 0) step <=   1105; else step = step + 1;/* endIfGe*/    end
         256 : begin if (intermediateValue != 0) step <=   1099; else step = step + 1;/* endIfNe*/    end
         257 : begin step <=   1105; /* end */ end
         258 : begin step <= 1089; /* start */ end
         259 : begin step <=   1205; /* end */ end
         260 : begin if (intermediateValue >= 0) step <=   1146; else step = step + 1;/* endIfGe*/    end
         261 : begin if (intermediateValue >  0) step <=   1140; else step = step + 1;/* endIfGt*/    end
         262 : begin step <=   1146; /* end */ end
         263 : begin step <= 1130; /* start */ end
         264 : begin if (intermediateValue == 0) step <=   1195; else step = step + 1;/* endIfEq*/    end
         265 : begin if (intermediateValue >= 0) step <=   1182; else step = step + 1;/* endIfGe*/    end
         266 : begin if (intermediateValue != 0) step <=   1176; else step = step + 1;/* endIfNe*/    end
         267 : begin step <=   1182; /* end */ end
         268 : begin step <= 1166; /* start */ end
         269 : begin if (intermediateValue >= 0) step <=   1204; else step = step + 1;/* endIfGe*/    end
         270 : begin step <= 1119; /* start */ end
         271 : begin if (intermediateValue == 0) step <=   1227; else step = step + 1;/* endIfEq*/    end
         272 : begin if (intermediateValue <  0) step <=   1224; else step = step + 1;/* endIfLt*/    end
         273 : begin step <=   1303; /* end */ end
         274 : begin if (intermediateValue >  0) step <=   1301; else step = step + 1;/* endIfGt*/    end
         275 : begin if (intermediateValue >= 0) step <=   1263; else step = step + 1;/* endIfGe*/    end
         276 : begin if (intermediateValue >  0) step <=   1257; else step = step + 1;/* endIfGt*/    end
         277 : begin step <=   1263; /* end */ end
         278 : begin step <= 1247; /* start */ end
         279 : begin if (intermediateValue == 0) step <=   1291; else step = step + 1;/* endIfEq*/    end
         280 : begin step <= 1278; /* start */ end
         281 : begin memory[249]/*merge_Key*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         282 : begin if (intermediateValue >  0) step <=   1936; else step = step + 1;/* endIfGt*/    end
         283 : begin memory[3] <= 0; /* clear 1 */ step <= step + 1; end
         284 : begin memory[279]/*mergeRoot_nP*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         285 : begin intermediateValue <= memory[279]/*mergeRoot_nP*/; /* get 1 */ step <= step + 1; end
         286 : begin intermediateValue <= 1 <  intermediateValue ? -1 : 1 == intermediateValue ?  0 : +1; /* compare 1 */ step <= step + 1; end
         287 : begin memory[276]/*mergeRoot_l*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         288 : begin memory[282]/*mergeRoot_r*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         289 : begin memory[141]/*hasLeavesForChildren*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         290 : begin intermediateValue <= memory[25+memory[141]/*hasLeavesForChildren*/*4+memory[0]]/*data[0,hasLeavesForChildren]*/; /* get 3 */ step <= step + 1; end
         291 : begin intermediateValue <= memory[141]/*hasLeavesForChildren*/; /* get 1 */ step <= step + 1; end
         292 : begin if (intermediateValue == 0) step <=   1570; else step = step + 1;/* endIfEq*/    end
         293 : begin intermediateValue <= memory[276]/*mergeRoot_l*/; /* get 1 */ step <= step + 1; end
         294 : begin memory[277]/*mergeRoot_nl*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         295 : begin intermediateValue <= memory[282]/*mergeRoot_r*/; /* get 1 */ step <= step + 1; end
         296 : begin memory[280]/*mergeRoot_nr*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         297 : begin intermediateValue <= memory[277]/*mergeRoot_nl*/; /* get 1 */ step <= step + 1; end
         298 : begin memory[278]/*mergeRoot_nlr*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         299 : begin intermediateValue <= memory[280]/*mergeRoot_nr*/ + memory[278]/*mergeRoot_nlr*/; /* add2 */ step <= step + 1; end
         300 : begin intermediateValue <= memory[278]/*mergeRoot_nlr*/; /* get 1 */ step <= step + 1; end
         301 : begin intermediateValue <= 0 <  intermediateValue ? -1 : 0 == intermediateValue ?  0 : +1; /* compare 1 */ step <= step + 1; end
         302 : begin if (intermediateValue <= 0) step <=   1453; else step = step + 1;/* endIfLe*/    end
         303 : begin if (intermediateValue >= 0) step <=   1398; else step = step + 1;/* endIfGe*/    end
         304 : begin step <= 1385; /* start */ end
         305 : begin if (intermediateValue >= 0) step <=   1439; else step = step + 1;/* endIfGe*/    end
         306 : begin step <= 1426; /* start */ end
         307 : begin intermediateValue <= memory[280]/*mergeRoot_nr*/; /* get 1 */ step <= step + 1; end
         308 : begin if (intermediateValue <= 0) step <=   1535; else step = step + 1;/* endIfLe*/    end
         309 : begin if (intermediateValue >= 0) step <=   1480; else step = step + 1;/* endIfGe*/    end
         310 : begin step <= 1467; /* start */ end
         311 : begin if (intermediateValue >= 0) step <=   1521; else step = step + 1;/* endIfGe*/    end
         312 : begin step <= 1508; /* start */ end
         313 : begin memory[120+memory[276]/*mergeRoot_l*/]/*free[mergeRoot_l]*/ <= -1; /* set 2 */ step <= step + 1; end
         314 : begin memory[145+memory[276]/*mergeRoot_l*/]/*isLeaf[mergeRoot_l]*/ <= -1; /* set 2 */ step <= step + 1; end
         315 : begin memory[5+memory[276]/*mergeRoot_l*/]/*current_size[mergeRoot_l]*/ <= -1; /* set 2 */ step <= step + 1; end
         316 : begin memory[166] <= -1; /* clear 2 */ step <= step + 1; end
         317 : begin memory[167] <= -1; /* clear 2 */ step <= step + 1; end
         318 : begin memory[168] <= -1; /* clear 2 */ step <= step + 1; end
         319 : begin memory[169] <= -1; /* clear 2 */ step <= step + 1; end
         320 : begin memory[25] <= -1; /* clear 2 */ step <= step + 1; end
         321 : begin memory[26] <= -1; /* clear 2 */ step <= step + 1; end
         322 : begin memory[27] <= -1; /* clear 2 */ step <= step + 1; end
         323 : begin memory[28] <= -1; /* clear 2 */ step <= step + 1; end
         324 : begin memory[120+memory[276]/*mergeRoot_l*/]/*free[mergeRoot_l]*/ <= intermediateValue; /* set 2 */ step <= step + 1; end
         325 : begin memory[120+memory[282]/*mergeRoot_r*/]/*free[mergeRoot_r]*/ <= -1; /* set 2 */ step <= step + 1; end
         326 : begin memory[145+memory[282]/*mergeRoot_r*/]/*isLeaf[mergeRoot_r]*/ <= -1; /* set 2 */ step <= step + 1; end
         327 : begin memory[5+memory[282]/*mergeRoot_r*/]/*current_size[mergeRoot_r]*/ <= -1; /* set 2 */ step <= step + 1; end
         328 : begin memory[120+memory[282]/*mergeRoot_r*/]/*free[mergeRoot_r]*/ <= intermediateValue; /* set 2 */ step <= step + 1; end
         329 : begin memory[281]/*mergeRoot_pkn*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         330 : begin if (intermediateValue <= 0) step <=   1733; else step = step + 1;/* endIfLe*/    end
         331 : begin if (intermediateValue >= 0) step <=   1637; else step = step + 1;/* endIfGe*/    end
         332 : begin step <= 1624; /* start */ end
         333 : begin if (intermediateValue >= 0) step <=   1678; else step = step + 1;/* endIfGe*/    end
         334 : begin step <= 1665; /* start */ end
         335 : begin if (intermediateValue >= 0) step <=   1719; else step = step + 1;/* endIfGe*/    end
         336 : begin step <= 1706; /* start */ end
         337 : begin intermediateValue <= memory[281]/*mergeRoot_pkn*/; /* get 1 */ step <= step + 1; end
         338 : begin if (intermediateValue <= 0) step <=   1880; else step = step + 1;/* endIfLe*/    end
         339 : begin if (intermediateValue >= 0) step <=   1784; else step = step + 1;/* endIfGe*/    end
         340 : begin step <= 1771; /* start */ end
         341 : begin if (intermediateValue >= 0) step <=   1825; else step = step + 1;/* endIfGe*/    end
         342 : begin step <= 1812; /* start */ end
         343 : begin if (intermediateValue >= 0) step <=   1866; else step = step + 1;/* endIfGe*/    end
         344 : begin step <= 1853; /* start */ end
         345 : begin memory[261] <= 0; /* clear 1 */ step <= step + 1; end
         346 : begin memory[261]/*merge_loop*/ <= 0; /* set 1 */ step <= step + 1; end
         347 : begin if (intermediateValue >  0) step <=   2868; else step = step + 1;/* endIfGt*/    end
         348 : begin memory[247]/*merge_indexLimit*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         349 : begin intermediateValue <= memory[247]/*merge_indexLimit*/; /* get 1 */ step <= step + 1; end
         350 : begin memory[248]/*merge_indices*/ <= 0; /* set 1 */ step <= step + 1; end
         351 : begin intermediateValue <= memory[248]/*merge_indices*/ < memory[247]/*merge_indexLimit*/ ? -1 : memory[248]/*merge_indices*/ == memory[247]/*merge_indexLimit*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
         352 : begin if (intermediateValue >= 0) step <=   2827; else step = step + 1;/* endIfGe*/    end
         353 : begin memory[256]/*mergeLeftSibling_parent*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         354 : begin intermediateValue <= memory[248]/*merge_indices*/; /* get 1 */ step <= step + 1; end
         355 : begin memory[251]/*mergeLeftSibling_index*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         356 : begin memory[260] <= 0; /* clear 1 */ step <= step + 1; end
         357 : begin intermediateValue <= memory[251]/*mergeLeftSibling_index*/; /* get 1 */ step <= step + 1; end
         358 : begin if (intermediateValue == 0) step <=   2395; else step = step + 1;/* endIfEq*/    end
         359 : begin intermediateValue <= memory[256]/*mergeLeftSibling_parent*/; /* get 1 */ step <= step + 1; end
         360 : begin memory[250]/*mergeLeftSibling_bs*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         361 : begin intermediateValue <= memory[251]/*mergeLeftSibling_index*/ < memory[250]/*mergeLeftSibling_bs*/ ? -1 : memory[251]/*mergeLeftSibling_index*/ == memory[250]/*mergeLeftSibling_bs*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
         362 : begin if (intermediateValue >= 0) step <=   2395; else step = step + 1;/* endIfGe*/    end
         363 : begin memory[252]/*mergeLeftSibling_l*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         364 : begin memory[257]/*mergeLeftSibling_r*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         365 : begin if (intermediateValue == 0) step <=   2113; else step = step + 1;/* endIfEq*/    end
         366 : begin intermediateValue <= memory[252]/*mergeLeftSibling_l*/; /* get 1 */ step <= step + 1; end
         367 : begin memory[253]/*mergeLeftSibling_nl*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         368 : begin intermediateValue <= memory[257]/*mergeLeftSibling_r*/; /* get 1 */ step <= step + 1; end
         369 : begin memory[255]/*mergeLeftSibling_nr*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         370 : begin intermediateValue <= memory[253]/*mergeLeftSibling_nl*/; /* get 1 */ step <= step + 1; end
         371 : begin memory[254]/*mergeLeftSibling_nlr*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         372 : begin intermediateValue <= memory[255]/*mergeLeftSibling_nr*/ + memory[254]/*mergeLeftSibling_nlr*/; /* add2 */ step <= step + 1; end
         373 : begin intermediateValue <= memory[254]/*mergeLeftSibling_nlr*/; /* get 1 */ step <= step + 1; end
         374 : begin intermediateValue <= memory[5+memory[252]/*mergeLeftSibling_l*/]/*current_size[mergeLeftSibling_l]*/; /* get 2 */ step <= step + 1; end
         375 : begin memory[258]/*mergeLeftSibling_size*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         376 : begin intermediateValue <= memory[258]/*mergeLeftSibling_size*/; /* get 1 */ step <= step + 1; end
         377 : begin if (intermediateValue <= 0) step <=   2113; else step = step + 1;/* endIfLe*/    end
         378 : begin memory[349]/*stuckUnshift_i*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         379 : begin intermediateValue <= memory[349]/*stuckUnshift_i*/; /* get 1 */ step <= step + 1; end
         380 : begin if (intermediateValue <= 0) step <=   2064; else step = step + 1;/* endIfLe*/    end
         381 : begin memory[350]/*stuckUnshift_I*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         382 : begin intermediateValue <= memory[350]/*stuckUnshift_I*/; /* get 1 */ step <= step + 1; end
         383 : begin intermediateValue <= memory[166+memory[348]/*stuck*/*4+memory[350]/*stuckUnshift_I*/]/*keys[stuckUnshift_I,stuck]*/; /* get 3 */ step <= step + 1; end
         384 : begin memory[166+memory[348]/*stuck*/*4+memory[349]/*stuckUnshift_i*/]/*keys[stuckUnshift_i,stuck]*/ <= intermediateValue; /* set 3 */ step <= step + 1; end
         385 : begin intermediateValue <= memory[25+memory[348]/*stuck*/*4+memory[350]/*stuckUnshift_I*/]/*data[stuckUnshift_I,stuck]*/; /* get 3 */ step <= step + 1; end
         386 : begin memory[25+memory[348]/*stuck*/*4+memory[349]/*stuckUnshift_i*/]/*data[stuckUnshift_i,stuck]*/ <= intermediateValue; /* set 3 */ step <= step + 1; end
         387 : begin step <= 2049; /* start */ end
         388 : begin if (intermediateValue <= 0) step <=   2105; else step = step + 1;/* endIfLe*/    end
         389 : begin step <= 2090; /* start */ end
         390 : begin if (intermediateValue >  0) step <=   2342; else step = step + 1;/* endIfGt*/    end
         391 : begin if (intermediateValue >  0) step <=   2395; else step = step + 1;/* endIfGt*/    end
         392 : begin memory[259]/*mergeLeftSibling_t*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         393 : begin intermediateValue <= memory[259]/*mergeLeftSibling_t*/; /* get 1 */ step <= step + 1; end
         394 : begin if (intermediateValue <= 0) step <=   2188; else step = step + 1;/* endIfLe*/    end
         395 : begin step <= 2173; /* start */ end
         396 : begin if (intermediateValue <= 0) step <=   2342; else step = step + 1;/* endIfLe*/    end
         397 : begin if (intermediateValue <= 0) step <=   2252; else step = step + 1;/* endIfLe*/    end
         398 : begin step <= 2237; /* start */ end
         399 : begin if (intermediateValue <= 0) step <=   2293; else step = step + 1;/* endIfLe*/    end
         400 : begin step <= 2278; /* start */ end
         401 : begin if (intermediateValue <= 0) step <=   2334; else step = step + 1;/* endIfLe*/    end
         402 : begin step <= 2319; /* start */ end
         403 : begin memory[120+memory[252]/*mergeLeftSibling_l*/]/*free[mergeLeftSibling_l]*/ <= -1; /* set 2 */ step <= step + 1; end
         404 : begin memory[145+memory[252]/*mergeLeftSibling_l*/]/*isLeaf[mergeLeftSibling_l]*/ <= -1; /* set 2 */ step <= step + 1; end
         405 : begin memory[5+memory[252]/*mergeLeftSibling_l*/]/*current_size[mergeLeftSibling_l]*/ <= -1; /* set 2 */ step <= step + 1; end
         406 : begin memory[120+memory[252]/*mergeLeftSibling_l*/]/*free[mergeLeftSibling_l]*/ <= intermediateValue; /* set 2 */ step <= step + 1; end
         407 : begin memory[343]/*stuckRemoveElementAt_N*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         408 : begin memory[342]/*stuckRemoveElementAt_i*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         409 : begin intermediateValue <= memory[342]/*stuckRemoveElementAt_i*/; /* get 1 */ step <= step + 1; end
         410 : begin memory[341]/*stuckRemoveElementAt_I*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         411 : begin intermediateValue <= memory[341]/*stuckRemoveElementAt_I*/; /* get 1 */ step <= step + 1; end
         412 : begin intermediateValue <= memory[341]/*stuckRemoveElementAt_I*/ < memory[343]/*stuckRemoveElementAt_N*/ ? -1 : memory[341]/*stuckRemoveElementAt_I*/ == memory[343]/*stuckRemoveElementAt_N*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
         413 : begin if (intermediateValue == 0) step <=   2391; else step = step + 1;/* endIfEq*/    end
         414 : begin intermediateValue <= memory[166+memory[348]/*stuck*/*4+memory[341]/*stuckRemoveElementAt_I*/]/*keys[stuckRemoveElementAt_I,stuck]*/; /* get 3 */ step <= step + 1; end
         415 : begin memory[166+memory[348]/*stuck*/*4+memory[342]/*stuckRemoveElementAt_i*/]/*keys[stuckRemoveElementAt_i,stuck]*/ <= intermediateValue; /* set 3 */ step <= step + 1; end
         416 : begin intermediateValue <= memory[25+memory[348]/*stuck*/*4+memory[341]/*stuckRemoveElementAt_I*/]/*data[stuckRemoveElementAt_I,stuck]*/; /* get 3 */ step <= step + 1; end
         417 : begin memory[25+memory[348]/*stuck*/*4+memory[342]/*stuckRemoveElementAt_i*/]/*data[stuckRemoveElementAt_i,stuck]*/ <= intermediateValue; /* set 3 */ step <= step + 1; end
         418 : begin step <= 2378; /* start */ end
         419 : begin memory[260] <= 1; /* clear 1 */ step <= step + 1; end
         420 : begin intermediateValue <= memory[260]/*mergeLeftSibling*/; /* get 1 */ step <= step + 1; end
         421 : begin if (intermediateValue == 0) step <=   2400; else step = step + 1;/* endIfEq*/    end
         422 : begin memory[248]/*merge_indices*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         423 : begin memory[270]/*mergeRightSibling_parent*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         424 : begin memory[264]/*mergeRightSibling_index*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         425 : begin memory[275] <= 0; /* clear 1 */ step <= step + 1; end
         426 : begin intermediateValue <= memory[5+memory[270]/*mergeRightSibling_parent*/]/*current_size[mergeRightSibling_parent]*/; /* get 2 */ step <= step + 1; end
         427 : begin memory[262]/*mergeRightSibling_bs*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         428 : begin intermediateValue <= memory[262]/*mergeRightSibling_bs*/; /* get 1 */ step <= step + 1; end
         429 : begin intermediateValue <= memory[264]/*mergeRightSibling_index*/ < memory[262]/*mergeRightSibling_bs*/ ? -1 : memory[264]/*mergeRightSibling_index*/ == memory[262]/*mergeRightSibling_bs*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
         430 : begin if (intermediateValue >= 0) step <=   2823; else step = step + 1;/* endIfGe*/    end
         431 : begin intermediateValue <= memory[270]/*mergeRightSibling_parent*/; /* get 1 */ step <= step + 1; end
         432 : begin intermediateValue <= memory[264]/*mergeRightSibling_index*/; /* get 1 */ step <= step + 1; end
         433 : begin memory[266]/*mergeRightSibling_l*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         434 : begin memory[272]/*mergeRightSibling_r*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         435 : begin if (intermediateValue == 0) step <=   2546; else step = step + 1;/* endIfEq*/    end
         436 : begin intermediateValue <= memory[266]/*mergeRightSibling_l*/; /* get 1 */ step <= step + 1; end
         437 : begin memory[267]/*mergeRightSibling_nl*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         438 : begin intermediateValue <= memory[272]/*mergeRightSibling_r*/; /* get 1 */ step <= step + 1; end
         439 : begin memory[269]/*mergeRightSibling_nr*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         440 : begin intermediateValue <= memory[267]/*mergeRightSibling_nl*/; /* get 1 */ step <= step + 1; end
         441 : begin memory[268]/*mergeRightSibling_nlr*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         442 : begin intermediateValue <= memory[269]/*mergeRightSibling_nr*/ + memory[268]/*mergeRightSibling_nlr*/; /* add2 */ step <= step + 1; end
         443 : begin intermediateValue <= memory[268]/*mergeRightSibling_nlr*/; /* get 1 */ step <= step + 1; end
         444 : begin if (intermediateValue >  0) step <=   2823; else step = step + 1;/* endIfGt*/    end
         445 : begin intermediateValue <= memory[5+memory[272]/*mergeRightSibling_r*/]/*current_size[mergeRightSibling_r]*/; /* get 2 */ step <= step + 1; end
         446 : begin memory[273]/*mergeRightSibling_size*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         447 : begin intermediateValue <= memory[273]/*mergeRightSibling_size*/; /* get 1 */ step <= step + 1; end
         448 : begin if (intermediateValue <= 0) step <=   2546; else step = step + 1;/* endIfLe*/    end
         449 : begin if (intermediateValue >= 0) step <=   2491; else step = step + 1;/* endIfGe*/    end
         450 : begin step <= 2478; /* start */ end
         451 : begin if (intermediateValue >= 0) step <=   2532; else step = step + 1;/* endIfGe*/    end
         452 : begin step <= 2519; /* start */ end
         453 : begin if (intermediateValue >  0) step <=   2740; else step = step + 1;/* endIfGt*/    end
         454 : begin memory[265]/*mergeRightSibling_ld*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         455 : begin intermediateValue <= memory[265]/*mergeRightSibling_ld*/; /* get 1 */ step <= step + 1; end
         456 : begin if (intermediateValue <  0) step <=   2612; else step = step + 1;/* endIfLt*/    end
         457 : begin intermediateValue <= memory[269]/*mergeRightSibling_nr*/; /* get 1 */ step <= step + 1; end
         458 : begin if (intermediateValue <= 0) step <=   2740; else step = step + 1;/* endIfLe*/    end
         459 : begin if (intermediateValue >= 0) step <=   2644; else step = step + 1;/* endIfGe*/    end
         460 : begin step <= 2631; /* start */ end
         461 : begin if (intermediateValue >= 0) step <=   2685; else step = step + 1;/* endIfGe*/    end
         462 : begin step <= 2672; /* start */ end
         463 : begin if (intermediateValue >= 0) step <=   2726; else step = step + 1;/* endIfGe*/    end
         464 : begin step <= 2713; /* start */ end
         465 : begin memory[120+memory[272]/*mergeRightSibling_r*/]/*free[mergeRightSibling_r]*/ <= -1; /* set 2 */ step <= step + 1; end
         466 : begin memory[145+memory[272]/*mergeRightSibling_r*/]/*isLeaf[mergeRightSibling_r]*/ <= -1; /* set 2 */ step <= step + 1; end
         467 : begin memory[5+memory[272]/*mergeRightSibling_r*/]/*current_size[mergeRightSibling_r]*/ <= -1; /* set 2 */ step <= step + 1; end
         468 : begin memory[120+memory[272]/*mergeRightSibling_r*/]/*free[mergeRightSibling_r]*/ <= intermediateValue; /* set 2 */ step <= step + 1; end
         469 : begin memory[271]/*mergeRightSibling_pk*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         470 : begin intermediateValue <= memory[271]/*mergeRightSibling_pk*/; /* get 1 */ step <= step + 1; end
         471 : begin if (intermediateValue <  0) step <=   2788; else step = step + 1;/* endIfLt*/    end
         472 : begin if (intermediateValue == 0) step <=   2819; else step = step + 1;/* endIfEq*/    end
         473 : begin step <= 2806; /* start */ end
         474 : begin memory[275] <= 1; /* clear 1 */ step <= step + 1; end
         475 : begin step <= 1959; /* start */ end
         476 : begin intermediateValue <= memory[249]/*merge_Key*/; /* get 1 */ step <= step + 1; end
         477 : begin if (intermediateValue >= 0) step <=   2854; else step = step + 1;/* endIfGe*/    end
         478 : begin if (intermediateValue >  0) step <=   2848; else step = step + 1;/* endIfGt*/    end
         479 : begin step <=   2854; /* end */ end
         480 : begin step <= 2838; /* start */ end
         481 : begin intermediateValue <= memory[261]/*merge_loop*/; /* get 1 */ step <= step + 1; end
         482 : begin memory[261]/*merge_loop*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         483 : begin if (intermediateValue >= 0) step <=   2867; else step = step + 1;/* endIfGe*/    end
         484 : begin step <= 1940; /* start */ end
         485 : begin step <=   3073; /* end */ end
         486 : begin if (intermediateValue == 0) step <=   3061; else step = step + 1;/* endIfEq*/    end
         487 : begin memory[297]/*splitBranch_node*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         488 : begin memory[298]/*splitBranch_parent*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         489 : begin memory[295]/*splitBranch_index*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         490 : begin memory[296]/*splitBranch_l*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         491 : begin intermediateValue <= memory[296]/*splitBranch_l*/; /* get 1 */ step <= step + 1; end
         492 : begin if (intermediateValue >  0) step <=   2895; else step = step + 1;/* endIfGt*/    end
         493 : begin intermediateValue <= memory[120+memory[296]/*splitBranch_l*/]/*free[splitBranch_l]*/; /* get 2 */ step <= step + 1; end
         494 : begin memory[120+memory[296]/*splitBranch_l*/]/*free[splitBranch_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         495 : begin memory[145+memory[296]/*splitBranch_l*/]/*isLeaf[splitBranch_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         496 : begin memory[5+memory[296]/*splitBranch_l*/]/*current_size[splitBranch_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         497 : begin intermediateValue <= memory[297]/*splitBranch_node*/; /* get 1 */ step <= step + 1; end
         498 : begin if (intermediateValue >= 0) step <=   2935; else step = step + 1;/* endIfGe*/    end
         499 : begin step <= 2922; /* start */ end
         500 : begin if (intermediateValue >= 0) step <=   2973; else step = step + 1;/* endIfGe*/    end
         501 : begin step <= 2960; /* start */ end
         502 : begin memory[299]/*splitBranch_rk*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         503 : begin intermediateValue <= memory[298]/*splitBranch_parent*/; /* get 1 */ step <= step + 1; end
         504 : begin intermediateValue <= memory[299]/*splitBranch_rk*/; /* get 1 */ step <= step + 1; end
         505 : begin intermediateValue <= memory[295]/*splitBranch_index*/; /* get 1 */ step <= step + 1; end
         506 : begin if (intermediateValue == 0) step <=   3021; else step = step + 1;/* endIfEq*/    end
         507 : begin step <= 3008; /* start */ end
         508 : begin if (intermediateValue >= 0) step <=   3055; else step = step + 1;/* endIfGe*/    end
         509 : begin if (intermediateValue >  0) step <=   3049; else step = step + 1;/* endIfGt*/    end
         510 : begin step <=   3055; /* end */ end
         511 : begin step <= 3039; /* start */ end
         512 : begin if (intermediateValue >  0) step <=   3065; else step = step + 1;/* endIfGt*/    end
         513 : begin intermediateValue <= memory[286]/*put_loop*/; /* get 1 */ step <= step + 1; end
         514 : begin memory[286]/*put_loop*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         515 : begin if (intermediateValue >  0) step <=   3072; else step = step + 1;/* endIfGt*/    end
         516 : begin step <= 906; /* start */ end

        default: stopped <= 1;
      endcase
      steps    <= steps + 1;
    end // Execute
  end // Always
endmodule
