//-----------------------------------------------------------------------------
// Generic cpu
// Philip R Brenan at appaapps dot com, Appa Apps Ltd Inc., 2025-01-07
//------------------------------------------------------------------------------
`timescale 10ps/1ps
(* keep_hierarchy = "yes" *)
module put_wide(reset, stop, clock, Key, Data, data, found);                    // Database on a chip
  input                      reset;                                             // Restart the program run sequence when this goes high
  input                      clock;                                             // Program counter clock
  input [16-1:0]  Key;                                             // Input key
  input [16-1:0] Data;                                             // Input data
  output                      stop;                                             // Program has stopped when this goes high
  output[16-1:0] data;                                             // Output data
  output                     found;                                             // Whether the key was found on put, find delete

  integer step;
  integer steps;
  integer stopped;
  integer intermediateValue;
  reg [16-1:0] memory [499-1: 0]; /* declareVerilogMemory */
  reg [10-1: 0] opCodes[5868 : 0];

  assign stop  = stopped > 0 ? 1 : 0;
  assign found = memory[184];  // found
  assign data  = memory[183];   // data

  always @ (posedge clock) begin                                                // Execute next step in program
    if (reset) begin                                                            // Reset
      step     <= 0;
      steps    <= 0;
      stopped  <= 0;
      begin /* initilizeVerilogMemory */
        integer i;
        for (i = 0; i < 499; i = i + 1) begin
          memory[i] <= 0;
        end
      end
      memory[ 195] <=    1; /* freeChainHead */
      memory[ 197] <=    2; /* free[1] */
      memory[ 198] <=    3; /* free[2] */
      memory[ 199] <=    4; /* free[3] */
      memory[ 200] <=    5; /* free[4] */
      memory[ 201] <=    6; /* free[5] */
      memory[ 202] <=    7; /* free[6] */
      memory[ 203] <=    8; /* free[7] */
      memory[ 204] <=    9; /* free[8] */
      memory[ 205] <=   10; /* free[9] */
      memory[ 206] <=   11; /* free[10] */
      memory[ 207] <=   12; /* free[11] */
      memory[ 208] <=   13; /* free[12] */
      memory[ 209] <=   14; /* free[13] */
      memory[ 210] <=   15; /* free[14] */
      memory[ 217] <=    1; /* isLeaf[0] */

      opCodes[0] <= 0;
      opCodes[1412] <= 0;
      opCodes[1933] <= 0;
      opCodes[5826] <= 0;
      opCodes[1] <= 1;
      opCodes[2] <= 2;
      opCodes[3] <= 3;
      opCodes[4] <= 4;
      opCodes[137] <= 4;
      opCodes[169] <= 4;
      opCodes[193] <= 4;
      opCodes[1178] <= 4;
      opCodes[1311] <= 4;
      opCodes[1343] <= 4;
      opCodes[1367] <= 4;
      opCodes[1706] <= 4;
      opCodes[1839] <= 4;
      opCodes[1871] <= 4;
      opCodes[1895] <= 4;
      opCodes[5] <= 5;
      opCodes[1179] <= 5;
      opCodes[1707] <= 5;
      opCodes[6] <= 6;
      opCodes[264] <= 6;
      opCodes[1180] <= 6;
      opCodes[1708] <= 6;
      opCodes[1935] <= 6;
      opCodes[7] <= 7;
      opCodes[265] <= 7;
      opCodes[1181] <= 7;
      opCodes[1709] <= 7;
      opCodes[1936] <= 7;
      opCodes[8] <= 8;
      opCodes[266] <= 8;
      opCodes[695] <= 8;
      opCodes[1182] <= 8;
      opCodes[1710] <= 8;
      opCodes[1937] <= 8;
      opCodes[9] <= 9;
      opCodes[10] <= 10;
      opCodes[1184] <= 10;
      opCodes[1712] <= 10;
      opCodes[1950] <= 10;
      opCodes[11] <= 11;
      opCodes[49] <= 11;
      opCodes[88] <= 11;
      opCodes[1185] <= 11;
      opCodes[1223] <= 11;
      opCodes[1262] <= 11;
      opCodes[1713] <= 11;
      opCodes[1751] <= 11;
      opCodes[1790] <= 11;
      opCodes[12] <= 12;
      opCodes[23] <= 12;
      opCodes[50] <= 12;
      opCodes[64] <= 12;
      opCodes[75] <= 12;
      opCodes[89] <= 12;
      opCodes[100] <= 12;
      opCodes[138] <= 12;
      opCodes[170] <= 12;
      opCodes[181] <= 12;
      opCodes[194] <= 12;
      opCodes[338] <= 12;
      opCodes[376] <= 12;
      opCodes[414] <= 12;
      opCodes[452] <= 12;
      opCodes[490] <= 12;
      opCodes[528] <= 12;
      opCodes[566] <= 12;
      opCodes[604] <= 12;
      opCodes[640] <= 12;
      opCodes[653] <= 12;
      opCodes[670] <= 12;
      opCodes[683] <= 12;
      opCodes[767] <= 12;
      opCodes[805] <= 12;
      opCodes[843] <= 12;
      opCodes[881] <= 12;
      opCodes[919] <= 12;
      opCodes[947] <= 12;
      opCodes[961] <= 12;
      opCodes[999] <= 12;
      opCodes[1037] <= 12;
      opCodes[1075] <= 12;
      opCodes[1113] <= 12;
      opCodes[1139] <= 12;
      opCodes[1153] <= 12;
      opCodes[1166] <= 12;
      opCodes[1186] <= 12;
      opCodes[1197] <= 12;
      opCodes[1224] <= 12;
      opCodes[1238] <= 12;
      opCodes[1249] <= 12;
      opCodes[1263] <= 12;
      opCodes[1274] <= 12;
      opCodes[1312] <= 12;
      opCodes[1344] <= 12;
      opCodes[1355] <= 12;
      opCodes[1368] <= 12;
      opCodes[1413] <= 12;
      opCodes[1427] <= 12;
      opCodes[1438] <= 12;
      opCodes[1492] <= 12;
      opCodes[1530] <= 12;
      opCodes[1568] <= 12;
      opCodes[1606] <= 12;
      opCodes[1644] <= 12;
      opCodes[1657] <= 12;
      opCodes[1672] <= 12;
      opCodes[1714] <= 12;
      opCodes[1725] <= 12;
      opCodes[1752] <= 12;
      opCodes[1766] <= 12;
      opCodes[1777] <= 12;
      opCodes[1791] <= 12;
      opCodes[1802] <= 12;
      opCodes[1840] <= 12;
      opCodes[1872] <= 12;
      opCodes[1883] <= 12;
      opCodes[1896] <= 12;
      opCodes[1953] <= 12;
      opCodes[1964] <= 12;
      opCodes[2008] <= 12;
      opCodes[2049] <= 12;
      opCodes[2090] <= 12;
      opCodes[2131] <= 12;
      opCodes[2172] <= 12;
      opCodes[2213] <= 12;
      opCodes[2254] <= 12;
      opCodes[2295] <= 12;
      opCodes[2336] <= 12;
      opCodes[2377] <= 12;
      opCodes[2418] <= 12;
      opCodes[2459] <= 12;
      opCodes[2500] <= 12;
      opCodes[2541] <= 12;
      opCodes[2582] <= 12;
      opCodes[2623] <= 12;
      opCodes[2750] <= 12;
      opCodes[2763] <= 12;
      opCodes[2804] <= 12;
      opCodes[2845] <= 12;
      opCodes[2886] <= 12;
      opCodes[2927] <= 12;
      opCodes[2968] <= 12;
      opCodes[3009] <= 12;
      opCodes[3050] <= 12;
      opCodes[3091] <= 12;
      opCodes[3133] <= 12;
      opCodes[3139] <= 12;
      opCodes[3156] <= 12;
      opCodes[3197] <= 12;
      opCodes[3238] <= 12;
      opCodes[3279] <= 12;
      opCodes[3320] <= 12;
      opCodes[3361] <= 12;
      opCodes[3402] <= 12;
      opCodes[3443] <= 12;
      opCodes[3484] <= 12;
      opCodes[3526] <= 12;
      opCodes[3532] <= 12;
      opCodes[3649] <= 12;
      opCodes[3657] <= 12;
      opCodes[3704] <= 12;
      opCodes[3745] <= 12;
      opCodes[3786] <= 12;
      opCodes[3827] <= 12;
      opCodes[3868] <= 12;
      opCodes[3909] <= 12;
      opCodes[3950] <= 12;
      opCodes[3991] <= 12;
      opCodes[4059] <= 12;
      opCodes[4072] <= 12;
      opCodes[4078] <= 12;
      opCodes[4112] <= 12;
      opCodes[4138] <= 12;
      opCodes[4179] <= 12;
      opCodes[4220] <= 12;
      opCodes[4261] <= 12;
      opCodes[4302] <= 12;
      opCodes[4343] <= 12;
      opCodes[4384] <= 12;
      opCodes[4425] <= 12;
      opCodes[4466] <= 12;
      opCodes[4541] <= 12;
      opCodes[4583] <= 12;
      opCodes[4594] <= 12;
      opCodes[4637] <= 12;
      opCodes[4678] <= 12;
      opCodes[4719] <= 12;
      opCodes[4760] <= 12;
      opCodes[4801] <= 12;
      opCodes[4842] <= 12;
      opCodes[4883] <= 12;
      opCodes[4924] <= 12;
      opCodes[4996] <= 12;
      opCodes[5006] <= 12;
      opCodes[5036] <= 12;
      opCodes[5077] <= 12;
      opCodes[5118] <= 12;
      opCodes[5159] <= 12;
      opCodes[5200] <= 12;
      opCodes[5241] <= 12;
      opCodes[5282] <= 12;
      opCodes[5323] <= 12;
      opCodes[5364] <= 12;
      opCodes[5434] <= 12;
      opCodes[5442] <= 12;
      opCodes[5446] <= 12;
      opCodes[5473] <= 12;
      opCodes[5500] <= 12;
      opCodes[5514] <= 12;
      opCodes[5525] <= 12;
      opCodes[5597] <= 12;
      opCodes[5635] <= 12;
      opCodes[5673] <= 12;
      opCodes[5711] <= 12;
      opCodes[5749] <= 12;
      opCodes[5777] <= 12;
      opCodes[5790] <= 12;
      opCodes[5827] <= 12;
      opCodes[5841] <= 12;
      opCodes[5852] <= 12;
      opCodes[13] <= 13;
      opCodes[51] <= 13;
      opCodes[90] <= 13;
      opCodes[171] <= 13;
      opCodes[1187] <= 13;
      opCodes[1225] <= 13;
      opCodes[1264] <= 13;
      opCodes[1345] <= 13;
      opCodes[1414] <= 13;
      opCodes[1715] <= 13;
      opCodes[1753] <= 13;
      opCodes[1792] <= 13;
      opCodes[1873] <= 13;
      opCodes[5501] <= 13;
      opCodes[5828] <= 13;
      opCodes[14] <= 14;
      opCodes[52] <= 14;
      opCodes[91] <= 14;
      opCodes[172] <= 14;
      opCodes[638] <= 14;
      opCodes[1188] <= 14;
      opCodes[1226] <= 14;
      opCodes[1265] <= 14;
      opCodes[1346] <= 14;
      opCodes[1415] <= 14;
      opCodes[1642] <= 14;
      opCodes[1716] <= 14;
      opCodes[1754] <= 14;
      opCodes[1793] <= 14;
      opCodes[1874] <= 14;
      opCodes[1951] <= 14;
      opCodes[2748] <= 14;
      opCodes[3726] <= 14;
      opCodes[3767] <= 14;
      opCodes[3808] <= 14;
      opCodes[3849] <= 14;
      opCodes[3890] <= 14;
      opCodes[3931] <= 14;
      opCodes[3972] <= 14;
      opCodes[4013] <= 14;
      opCodes[4096] <= 14;
      opCodes[4160] <= 14;
      opCodes[4201] <= 14;
      opCodes[4242] <= 14;
      opCodes[4283] <= 14;
      opCodes[4324] <= 14;
      opCodes[4365] <= 14;
      opCodes[4406] <= 14;
      opCodes[4447] <= 14;
      opCodes[4488] <= 14;
      opCodes[5502] <= 14;
      opCodes[5829] <= 14;
      opCodes[15] <= 15;
      opCodes[53] <= 15;
      opCodes[92] <= 15;
      opCodes[149] <= 15;
      opCodes[173] <= 15;
      opCodes[199] <= 15;
      opCodes[223] <= 15;
      opCodes[341] <= 15;
      opCodes[358] <= 15;
      opCodes[363] <= 15;
      opCodes[369] <= 15;
      opCodes[379] <= 15;
      opCodes[396] <= 15;
      opCodes[401] <= 15;
      opCodes[407] <= 15;
      opCodes[417] <= 15;
      opCodes[434] <= 15;
      opCodes[439] <= 15;
      opCodes[445] <= 15;
      opCodes[455] <= 15;
      opCodes[472] <= 15;
      opCodes[477] <= 15;
      opCodes[483] <= 15;
      opCodes[493] <= 15;
      opCodes[510] <= 15;
      opCodes[515] <= 15;
      opCodes[521] <= 15;
      opCodes[531] <= 15;
      opCodes[548] <= 15;
      opCodes[553] <= 15;
      opCodes[559] <= 15;
      opCodes[569] <= 15;
      opCodes[586] <= 15;
      opCodes[591] <= 15;
      opCodes[597] <= 15;
      opCodes[607] <= 15;
      opCodes[624] <= 15;
      opCodes[629] <= 15;
      opCodes[635] <= 15;
      opCodes[647] <= 15;
      opCodes[673] <= 15;
      opCodes[679] <= 15;
      opCodes[686] <= 15;
      opCodes[692] <= 15;
      opCodes[770] <= 15;
      opCodes[787] <= 15;
      opCodes[792] <= 15;
      opCodes[798] <= 15;
      opCodes[808] <= 15;
      opCodes[825] <= 15;
      opCodes[830] <= 15;
      opCodes[836] <= 15;
      opCodes[846] <= 15;
      opCodes[863] <= 15;
      opCodes[868] <= 15;
      opCodes[874] <= 15;
      opCodes[884] <= 15;
      opCodes[901] <= 15;
      opCodes[906] <= 15;
      opCodes[912] <= 15;
      opCodes[922] <= 15;
      opCodes[939] <= 15;
      opCodes[948] <= 15;
      opCodes[954] <= 15;
      opCodes[964] <= 15;
      opCodes[981] <= 15;
      opCodes[986] <= 15;
      opCodes[992] <= 15;
      opCodes[1002] <= 15;
      opCodes[1019] <= 15;
      opCodes[1024] <= 15;
      opCodes[1030] <= 15;
      opCodes[1040] <= 15;
      opCodes[1057] <= 15;
      opCodes[1062] <= 15;
      opCodes[1068] <= 15;
      opCodes[1078] <= 15;
      opCodes[1095] <= 15;
      opCodes[1100] <= 15;
      opCodes[1106] <= 15;
      opCodes[1116] <= 15;
      opCodes[1133] <= 15;
      opCodes[1140] <= 15;
      opCodes[1146] <= 15;
      opCodes[1156] <= 15;
      opCodes[1162] <= 15;
      opCodes[1169] <= 15;
      opCodes[1175] <= 15;
      opCodes[1189] <= 15;
      opCodes[1227] <= 15;
      opCodes[1266] <= 15;
      opCodes[1323] <= 15;
      opCodes[1347] <= 15;
      opCodes[1373] <= 15;
      opCodes[1397] <= 15;
      opCodes[1416] <= 15;
      opCodes[1495] <= 15;
      opCodes[1512] <= 15;
      opCodes[1517] <= 15;
      opCodes[1523] <= 15;
      opCodes[1533] <= 15;
      opCodes[1550] <= 15;
      opCodes[1555] <= 15;
      opCodes[1561] <= 15;
      opCodes[1571] <= 15;
      opCodes[1588] <= 15;
      opCodes[1593] <= 15;
      opCodes[1599] <= 15;
      opCodes[1609] <= 15;
      opCodes[1626] <= 15;
      opCodes[1631] <= 15;
      opCodes[1637] <= 15;
      opCodes[1651] <= 15;
      opCodes[1679] <= 15;
      opCodes[1703] <= 15;
      opCodes[1717] <= 15;
      opCodes[1755] <= 15;
      opCodes[1794] <= 15;
      opCodes[1851] <= 15;
      opCodes[1875] <= 15;
      opCodes[1901] <= 15;
      opCodes[1925] <= 15;
      opCodes[1958] <= 15;
      opCodes[2011] <= 15;
      opCodes[2028] <= 15;
      opCodes[2033] <= 15;
      opCodes[2039] <= 15;
      opCodes[2052] <= 15;
      opCodes[2069] <= 15;
      opCodes[2074] <= 15;
      opCodes[2080] <= 15;
      opCodes[2093] <= 15;
      opCodes[2110] <= 15;
      opCodes[2115] <= 15;
      opCodes[2121] <= 15;
      opCodes[2134] <= 15;
      opCodes[2151] <= 15;
      opCodes[2156] <= 15;
      opCodes[2162] <= 15;
      opCodes[2175] <= 15;
      opCodes[2192] <= 15;
      opCodes[2197] <= 15;
      opCodes[2203] <= 15;
      opCodes[2216] <= 15;
      opCodes[2233] <= 15;
      opCodes[2238] <= 15;
      opCodes[2244] <= 15;
      opCodes[2257] <= 15;
      opCodes[2274] <= 15;
      opCodes[2279] <= 15;
      opCodes[2285] <= 15;
      opCodes[2298] <= 15;
      opCodes[2315] <= 15;
      opCodes[2320] <= 15;
      opCodes[2326] <= 15;
      opCodes[2339] <= 15;
      opCodes[2356] <= 15;
      opCodes[2361] <= 15;
      opCodes[2367] <= 15;
      opCodes[2380] <= 15;
      opCodes[2397] <= 15;
      opCodes[2402] <= 15;
      opCodes[2408] <= 15;
      opCodes[2421] <= 15;
      opCodes[2438] <= 15;
      opCodes[2443] <= 15;
      opCodes[2449] <= 15;
      opCodes[2462] <= 15;
      opCodes[2479] <= 15;
      opCodes[2484] <= 15;
      opCodes[2490] <= 15;
      opCodes[2503] <= 15;
      opCodes[2520] <= 15;
      opCodes[2525] <= 15;
      opCodes[2531] <= 15;
      opCodes[2544] <= 15;
      opCodes[2561] <= 15;
      opCodes[2566] <= 15;
      opCodes[2572] <= 15;
      opCodes[2585] <= 15;
      opCodes[2602] <= 15;
      opCodes[2607] <= 15;
      opCodes[2613] <= 15;
      opCodes[2626] <= 15;
      opCodes[2643] <= 15;
      opCodes[2648] <= 15;
      opCodes[2654] <= 15;
      opCodes[2766] <= 15;
      opCodes[2783] <= 15;
      opCodes[2788] <= 15;
      opCodes[2794] <= 15;
      opCodes[2807] <= 15;
      opCodes[2824] <= 15;
      opCodes[2829] <= 15;
      opCodes[2835] <= 15;
      opCodes[2848] <= 15;
      opCodes[2865] <= 15;
      opCodes[2870] <= 15;
      opCodes[2876] <= 15;
      opCodes[2889] <= 15;
      opCodes[2906] <= 15;
      opCodes[2911] <= 15;
      opCodes[2917] <= 15;
      opCodes[2930] <= 15;
      opCodes[2947] <= 15;
      opCodes[2952] <= 15;
      opCodes[2958] <= 15;
      opCodes[2971] <= 15;
      opCodes[2988] <= 15;
      opCodes[2993] <= 15;
      opCodes[2999] <= 15;
      opCodes[3012] <= 15;
      opCodes[3029] <= 15;
      opCodes[3034] <= 15;
      opCodes[3040] <= 15;
      opCodes[3053] <= 15;
      opCodes[3070] <= 15;
      opCodes[3075] <= 15;
      opCodes[3081] <= 15;
      opCodes[3094] <= 15;
      opCodes[3111] <= 15;
      opCodes[3116] <= 15;
      opCodes[3122] <= 15;
      opCodes[3127] <= 15;
      opCodes[3140] <= 15;
      opCodes[3146] <= 15;
      opCodes[3159] <= 15;
      opCodes[3176] <= 15;
      opCodes[3181] <= 15;
      opCodes[3187] <= 15;
      opCodes[3200] <= 15;
      opCodes[3217] <= 15;
      opCodes[3222] <= 15;
      opCodes[3228] <= 15;
      opCodes[3241] <= 15;
      opCodes[3258] <= 15;
      opCodes[3263] <= 15;
      opCodes[3269] <= 15;
      opCodes[3282] <= 15;
      opCodes[3299] <= 15;
      opCodes[3304] <= 15;
      opCodes[3310] <= 15;
      opCodes[3323] <= 15;
      opCodes[3340] <= 15;
      opCodes[3345] <= 15;
      opCodes[3351] <= 15;
      opCodes[3364] <= 15;
      opCodes[3381] <= 15;
      opCodes[3386] <= 15;
      opCodes[3392] <= 15;
      opCodes[3405] <= 15;
      opCodes[3422] <= 15;
      opCodes[3427] <= 15;
      opCodes[3433] <= 15;
      opCodes[3446] <= 15;
      opCodes[3463] <= 15;
      opCodes[3468] <= 15;
      opCodes[3474] <= 15;
      opCodes[3487] <= 15;
      opCodes[3504] <= 15;
      opCodes[3509] <= 15;
      opCodes[3515] <= 15;
      opCodes[3520] <= 15;
      opCodes[3533] <= 15;
      opCodes[3539] <= 15;
      opCodes[3698] <= 15;
      opCodes[3701] <= 15;
      opCodes[3709] <= 15;
      opCodes[3731] <= 15;
      opCodes[3739] <= 15;
      opCodes[3742] <= 15;
      opCodes[3750] <= 15;
      opCodes[3772] <= 15;
      opCodes[3780] <= 15;
      opCodes[3783] <= 15;
      opCodes[3791] <= 15;
      opCodes[3813] <= 15;
      opCodes[3821] <= 15;
      opCodes[3824] <= 15;
      opCodes[3832] <= 15;
      opCodes[3854] <= 15;
      opCodes[3862] <= 15;
      opCodes[3865] <= 15;
      opCodes[3873] <= 15;
      opCodes[3895] <= 15;
      opCodes[3903] <= 15;
      opCodes[3906] <= 15;
      opCodes[3914] <= 15;
      opCodes[3936] <= 15;
      opCodes[3944] <= 15;
      opCodes[3947] <= 15;
      opCodes[3955] <= 15;
      opCodes[3977] <= 15;
      opCodes[3985] <= 15;
      opCodes[3988] <= 15;
      opCodes[3996] <= 15;
      opCodes[4018] <= 15;
      opCodes[4066] <= 15;
      opCodes[4079] <= 15;
      opCodes[4101] <= 15;
      opCodes[4106] <= 15;
      opCodes[4109] <= 15;
      opCodes[4132] <= 15;
      opCodes[4135] <= 15;
      opCodes[4143] <= 15;
      opCodes[4165] <= 15;
      opCodes[4173] <= 15;
      opCodes[4176] <= 15;
      opCodes[4184] <= 15;
      opCodes[4206] <= 15;
      opCodes[4214] <= 15;
      opCodes[4217] <= 15;
      opCodes[4225] <= 15;
      opCodes[4247] <= 15;
      opCodes[4255] <= 15;
      opCodes[4258] <= 15;
      opCodes[4266] <= 15;
      opCodes[4288] <= 15;
      opCodes[4296] <= 15;
      opCodes[4299] <= 15;
      opCodes[4307] <= 15;
      opCodes[4329] <= 15;
      opCodes[4337] <= 15;
      opCodes[4340] <= 15;
      opCodes[4348] <= 15;
      opCodes[4370] <= 15;
      opCodes[4378] <= 15;
      opCodes[4381] <= 15;
      opCodes[4389] <= 15;
      opCodes[4411] <= 15;
      opCodes[4419] <= 15;
      opCodes[4422] <= 15;
      opCodes[4430] <= 15;
      opCodes[4452] <= 15;
      opCodes[4460] <= 15;
      opCodes[4463] <= 15;
      opCodes[4471] <= 15;
      opCodes[4493] <= 15;
      opCodes[4531] <= 15;
      opCodes[4557] <= 15;
      opCodes[4640] <= 15;
      opCodes[4657] <= 15;
      opCodes[4662] <= 15;
      opCodes[4668] <= 15;
      opCodes[4681] <= 15;
      opCodes[4698] <= 15;
      opCodes[4703] <= 15;
      opCodes[4709] <= 15;
      opCodes[4722] <= 15;
      opCodes[4739] <= 15;
      opCodes[4744] <= 15;
      opCodes[4750] <= 15;
      opCodes[4763] <= 15;
      opCodes[4780] <= 15;
      opCodes[4785] <= 15;
      opCodes[4791] <= 15;
      opCodes[4804] <= 15;
      opCodes[4821] <= 15;
      opCodes[4826] <= 15;
      opCodes[4832] <= 15;
      opCodes[4845] <= 15;
      opCodes[4862] <= 15;
      opCodes[4867] <= 15;
      opCodes[4873] <= 15;
      opCodes[4886] <= 15;
      opCodes[4903] <= 15;
      opCodes[4908] <= 15;
      opCodes[4914] <= 15;
      opCodes[4927] <= 15;
      opCodes[4944] <= 15;
      opCodes[4949] <= 15;
      opCodes[4955] <= 15;
      opCodes[4990] <= 15;
      opCodes[5021] <= 15;
      opCodes[5039] <= 15;
      opCodes[5056] <= 15;
      opCodes[5061] <= 15;
      opCodes[5067] <= 15;
      opCodes[5080] <= 15;
      opCodes[5097] <= 15;
      opCodes[5102] <= 15;
      opCodes[5108] <= 15;
      opCodes[5121] <= 15;
      opCodes[5138] <= 15;
      opCodes[5143] <= 15;
      opCodes[5149] <= 15;
      opCodes[5162] <= 15;
      opCodes[5179] <= 15;
      opCodes[5184] <= 15;
      opCodes[5190] <= 15;
      opCodes[5203] <= 15;
      opCodes[5220] <= 15;
      opCodes[5225] <= 15;
      opCodes[5231] <= 15;
      opCodes[5244] <= 15;
      opCodes[5261] <= 15;
      opCodes[5266] <= 15;
      opCodes[5272] <= 15;
      opCodes[5285] <= 15;
      opCodes[5302] <= 15;
      opCodes[5307] <= 15;
      opCodes[5313] <= 15;
      opCodes[5326] <= 15;
      opCodes[5343] <= 15;
      opCodes[5348] <= 15;
      opCodes[5354] <= 15;
      opCodes[5367] <= 15;
      opCodes[5384] <= 15;
      opCodes[5389] <= 15;
      opCodes[5395] <= 15;
      opCodes[5455] <= 15;
      opCodes[5463] <= 15;
      opCodes[5489] <= 15;
      opCodes[5503] <= 15;
      opCodes[5600] <= 15;
      opCodes[5617] <= 15;
      opCodes[5622] <= 15;
      opCodes[5628] <= 15;
      opCodes[5638] <= 15;
      opCodes[5655] <= 15;
      opCodes[5660] <= 15;
      opCodes[5666] <= 15;
      opCodes[5676] <= 15;
      opCodes[5693] <= 15;
      opCodes[5698] <= 15;
      opCodes[5704] <= 15;
      opCodes[5714] <= 15;
      opCodes[5731] <= 15;
      opCodes[5736] <= 15;
      opCodes[5742] <= 15;
      opCodes[5752] <= 15;
      opCodes[5769] <= 15;
      opCodes[5778] <= 15;
      opCodes[5784] <= 15;
      opCodes[5797] <= 15;
      opCodes[5821] <= 15;
      opCodes[5830] <= 15;
      opCodes[16] <= 16;
      opCodes[54] <= 16;
      opCodes[57] <= 16;
      opCodes[93] <= 16;
      opCodes[174] <= 16;
      opCodes[1190] <= 16;
      opCodes[1228] <= 16;
      opCodes[1231] <= 16;
      opCodes[1267] <= 16;
      opCodes[1348] <= 16;
      opCodes[1417] <= 16;
      opCodes[1420] <= 16;
      opCodes[1718] <= 16;
      opCodes[1756] <= 16;
      opCodes[1759] <= 16;
      opCodes[1795] <= 16;
      opCodes[1876] <= 16;
      opCodes[5504] <= 16;
      opCodes[5507] <= 16;
      opCodes[5831] <= 16;
      opCodes[5834] <= 16;
      opCodes[17] <= 17;
      opCodes[30] <= 17;
      opCodes[58] <= 17;
      opCodes[71] <= 17;
      opCodes[94] <= 17;
      opCodes[107] <= 17;
      opCodes[175] <= 17;
      opCodes[188] <= 17;
      opCodes[1191] <= 17;
      opCodes[1204] <= 17;
      opCodes[1232] <= 17;
      opCodes[1245] <= 17;
      opCodes[1268] <= 17;
      opCodes[1281] <= 17;
      opCodes[1349] <= 17;
      opCodes[1362] <= 17;
      opCodes[1421] <= 17;
      opCodes[1434] <= 17;
      opCodes[1719] <= 17;
      opCodes[1732] <= 17;
      opCodes[1760] <= 17;
      opCodes[1773] <= 17;
      opCodes[1796] <= 17;
      opCodes[1809] <= 17;
      opCodes[1877] <= 17;
      opCodes[1890] <= 17;
      opCodes[5508] <= 17;
      opCodes[5521] <= 17;
      opCodes[5835] <= 17;
      opCodes[5848] <= 17;
      opCodes[18] <= 18;
      opCodes[31] <= 18;
      opCodes[19] <= 19;
      opCodes[60] <= 19;
      opCodes[96] <= 19;
      opCodes[177] <= 19;
      opCodes[1193] <= 19;
      opCodes[1234] <= 19;
      opCodes[1270] <= 19;
      opCodes[1351] <= 19;
      opCodes[1423] <= 19;
      opCodes[1721] <= 19;
      opCodes[1762] <= 19;
      opCodes[1798] <= 19;
      opCodes[1879] <= 19;
      opCodes[5510] <= 19;
      opCodes[5837] <= 19;
      opCodes[20] <= 20;
      opCodes[21] <= 21;
      opCodes[62] <= 21;
      opCodes[98] <= 21;
      opCodes[179] <= 21;
      opCodes[1195] <= 21;
      opCodes[1236] <= 21;
      opCodes[1272] <= 21;
      opCodes[1353] <= 21;
      opCodes[1425] <= 21;
      opCodes[1723] <= 21;
      opCodes[1764] <= 21;
      opCodes[1800] <= 21;
      opCodes[1881] <= 21;
      opCodes[5512] <= 21;
      opCodes[5839] <= 21;
      opCodes[22] <= 22;
      opCodes[63] <= 22;
      opCodes[74] <= 22;
      opCodes[99] <= 22;
      opCodes[180] <= 22;
      opCodes[337] <= 22;
      opCodes[375] <= 22;
      opCodes[413] <= 22;
      opCodes[451] <= 22;
      opCodes[489] <= 22;
      opCodes[527] <= 22;
      opCodes[565] <= 22;
      opCodes[603] <= 22;
      opCodes[639] <= 22;
      opCodes[652] <= 22;
      opCodes[766] <= 22;
      opCodes[804] <= 22;
      opCodes[842] <= 22;
      opCodes[880] <= 22;
      opCodes[918] <= 22;
      opCodes[960] <= 22;
      opCodes[998] <= 22;
      opCodes[1036] <= 22;
      opCodes[1074] <= 22;
      opCodes[1112] <= 22;
      opCodes[1196] <= 22;
      opCodes[1237] <= 22;
      opCodes[1248] <= 22;
      opCodes[1273] <= 22;
      opCodes[1354] <= 22;
      opCodes[1426] <= 22;
      opCodes[1437] <= 22;
      opCodes[1491] <= 22;
      opCodes[1529] <= 22;
      opCodes[1567] <= 22;
      opCodes[1605] <= 22;
      opCodes[1643] <= 22;
      opCodes[1656] <= 22;
      opCodes[1724] <= 22;
      opCodes[1765] <= 22;
      opCodes[1776] <= 22;
      opCodes[1801] <= 22;
      opCodes[1882] <= 22;
      opCodes[1952] <= 22;
      opCodes[1963] <= 22;
      opCodes[2007] <= 22;
      opCodes[2048] <= 22;
      opCodes[2089] <= 22;
      opCodes[2130] <= 22;
      opCodes[2171] <= 22;
      opCodes[2212] <= 22;
      opCodes[2253] <= 22;
      opCodes[2294] <= 22;
      opCodes[2335] <= 22;
      opCodes[2376] <= 22;
      opCodes[2417] <= 22;
      opCodes[2458] <= 22;
      opCodes[2499] <= 22;
      opCodes[2540] <= 22;
      opCodes[2581] <= 22;
      opCodes[2622] <= 22;
      opCodes[2749] <= 22;
      opCodes[2762] <= 22;
      opCodes[2803] <= 22;
      opCodes[2844] <= 22;
      opCodes[2885] <= 22;
      opCodes[2926] <= 22;
      opCodes[2967] <= 22;
      opCodes[3008] <= 22;
      opCodes[3049] <= 22;
      opCodes[3090] <= 22;
      opCodes[3132] <= 22;
      opCodes[3155] <= 22;
      opCodes[3196] <= 22;
      opCodes[3237] <= 22;
      opCodes[3278] <= 22;
      opCodes[3319] <= 22;
      opCodes[3360] <= 22;
      opCodes[3401] <= 22;
      opCodes[3442] <= 22;
      opCodes[3483] <= 22;
      opCodes[3525] <= 22;
      opCodes[3648] <= 22;
      opCodes[3656] <= 22;
      opCodes[3703] <= 22;
      opCodes[3744] <= 22;
      opCodes[3785] <= 22;
      opCodes[3826] <= 22;
      opCodes[3867] <= 22;
      opCodes[3908] <= 22;
      opCodes[3949] <= 22;
      opCodes[3990] <= 22;
      opCodes[4058] <= 22;
      opCodes[4071] <= 22;
      opCodes[4111] <= 22;
      opCodes[4137] <= 22;
      opCodes[4178] <= 22;
      opCodes[4219] <= 22;
      opCodes[4260] <= 22;
      opCodes[4301] <= 22;
      opCodes[4342] <= 22;
      opCodes[4383] <= 22;
      opCodes[4424] <= 22;
      opCodes[4465] <= 22;
      opCodes[4540] <= 22;
      opCodes[4582] <= 22;
      opCodes[4593] <= 22;
      opCodes[4636] <= 22;
      opCodes[4677] <= 22;
      opCodes[4718] <= 22;
      opCodes[4759] <= 22;
      opCodes[4800] <= 22;
      opCodes[4841] <= 22;
      opCodes[4882] <= 22;
      opCodes[4923] <= 22;
      opCodes[4995] <= 22;
      opCodes[5005] <= 22;
      opCodes[5035] <= 22;
      opCodes[5076] <= 22;
      opCodes[5117] <= 22;
      opCodes[5158] <= 22;
      opCodes[5199] <= 22;
      opCodes[5240] <= 22;
      opCodes[5281] <= 22;
      opCodes[5322] <= 22;
      opCodes[5363] <= 22;
      opCodes[5433] <= 22;
      opCodes[5441] <= 22;
      opCodes[5472] <= 22;
      opCodes[5513] <= 22;
      opCodes[5524] <= 22;
      opCodes[5596] <= 22;
      opCodes[5634] <= 22;
      opCodes[5672] <= 22;
      opCodes[5710] <= 22;
      opCodes[5748] <= 22;
      opCodes[5840] <= 22;
      opCodes[5851] <= 22;
      opCodes[24] <= 23;
      opCodes[65] <= 23;
      opCodes[76] <= 23;
      opCodes[101] <= 23;
      opCodes[182] <= 23;
      opCodes[339] <= 23;
      opCodes[377] <= 23;
      opCodes[415] <= 23;
      opCodes[453] <= 23;
      opCodes[491] <= 23;
      opCodes[529] <= 23;
      opCodes[567] <= 23;
      opCodes[605] <= 23;
      opCodes[641] <= 23;
      opCodes[654] <= 23;
      opCodes[768] <= 23;
      opCodes[806] <= 23;
      opCodes[844] <= 23;
      opCodes[882] <= 23;
      opCodes[920] <= 23;
      opCodes[962] <= 23;
      opCodes[1000] <= 23;
      opCodes[1038] <= 23;
      opCodes[1076] <= 23;
      opCodes[1114] <= 23;
      opCodes[1198] <= 23;
      opCodes[1239] <= 23;
      opCodes[1250] <= 23;
      opCodes[1275] <= 23;
      opCodes[1356] <= 23;
      opCodes[1428] <= 23;
      opCodes[1439] <= 23;
      opCodes[1493] <= 23;
      opCodes[1531] <= 23;
      opCodes[1569] <= 23;
      opCodes[1607] <= 23;
      opCodes[1645] <= 23;
      opCodes[1658] <= 23;
      opCodes[1726] <= 23;
      opCodes[1767] <= 23;
      opCodes[1778] <= 23;
      opCodes[1803] <= 23;
      opCodes[1884] <= 23;
      opCodes[1954] <= 23;
      opCodes[1965] <= 23;
      opCodes[2009] <= 23;
      opCodes[2050] <= 23;
      opCodes[2091] <= 23;
      opCodes[2132] <= 23;
      opCodes[2173] <= 23;
      opCodes[2214] <= 23;
      opCodes[2255] <= 23;
      opCodes[2296] <= 23;
      opCodes[2337] <= 23;
      opCodes[2378] <= 23;
      opCodes[2419] <= 23;
      opCodes[2460] <= 23;
      opCodes[2501] <= 23;
      opCodes[2542] <= 23;
      opCodes[2583] <= 23;
      opCodes[2624] <= 23;
      opCodes[2751] <= 23;
      opCodes[2764] <= 23;
      opCodes[2805] <= 23;
      opCodes[2846] <= 23;
      opCodes[2887] <= 23;
      opCodes[2928] <= 23;
      opCodes[2969] <= 23;
      opCodes[3010] <= 23;
      opCodes[3051] <= 23;
      opCodes[3092] <= 23;
      opCodes[3134] <= 23;
      opCodes[3157] <= 23;
      opCodes[3198] <= 23;
      opCodes[3239] <= 23;
      opCodes[3280] <= 23;
      opCodes[3321] <= 23;
      opCodes[3362] <= 23;
      opCodes[3403] <= 23;
      opCodes[3444] <= 23;
      opCodes[3485] <= 23;
      opCodes[3527] <= 23;
      opCodes[3650] <= 23;
      opCodes[3658] <= 23;
      opCodes[3705] <= 23;
      opCodes[3746] <= 23;
      opCodes[3787] <= 23;
      opCodes[3828] <= 23;
      opCodes[3869] <= 23;
      opCodes[3910] <= 23;
      opCodes[3951] <= 23;
      opCodes[3992] <= 23;
      opCodes[4060] <= 23;
      opCodes[4073] <= 23;
      opCodes[4113] <= 23;
      opCodes[4139] <= 23;
      opCodes[4180] <= 23;
      opCodes[4221] <= 23;
      opCodes[4262] <= 23;
      opCodes[4303] <= 23;
      opCodes[4344] <= 23;
      opCodes[4385] <= 23;
      opCodes[4426] <= 23;
      opCodes[4467] <= 23;
      opCodes[4542] <= 23;
      opCodes[4584] <= 23;
      opCodes[4595] <= 23;
      opCodes[4638] <= 23;
      opCodes[4679] <= 23;
      opCodes[4720] <= 23;
      opCodes[4761] <= 23;
      opCodes[4802] <= 23;
      opCodes[4843] <= 23;
      opCodes[4884] <= 23;
      opCodes[4925] <= 23;
      opCodes[4997] <= 23;
      opCodes[5007] <= 23;
      opCodes[5037] <= 23;
      opCodes[5078] <= 23;
      opCodes[5119] <= 23;
      opCodes[5160] <= 23;
      opCodes[5201] <= 23;
      opCodes[5242] <= 23;
      opCodes[5283] <= 23;
      opCodes[5324] <= 23;
      opCodes[5365] <= 23;
      opCodes[5435] <= 23;
      opCodes[5443] <= 23;
      opCodes[5474] <= 23;
      opCodes[5515] <= 23;
      opCodes[5526] <= 23;
      opCodes[5598] <= 23;
      opCodes[5636] <= 23;
      opCodes[5674] <= 23;
      opCodes[5712] <= 23;
      opCodes[5750] <= 23;
      opCodes[5842] <= 23;
      opCodes[5853] <= 23;
      opCodes[25] <= 24;
      opCodes[66] <= 24;
      opCodes[77] <= 24;
      opCodes[102] <= 24;
      opCodes[140] <= 24;
      opCodes[183] <= 24;
      opCodes[196] <= 24;
      opCodes[340] <= 24;
      opCodes[378] <= 24;
      opCodes[416] <= 24;
      opCodes[454] <= 24;
      opCodes[492] <= 24;
      opCodes[530] <= 24;
      opCodes[568] <= 24;
      opCodes[606] <= 24;
      opCodes[642] <= 24;
      opCodes[655] <= 24;
      opCodes[672] <= 24;
      opCodes[685] <= 24;
      opCodes[769] <= 24;
      opCodes[807] <= 24;
      opCodes[845] <= 24;
      opCodes[883] <= 24;
      opCodes[921] <= 24;
      opCodes[963] <= 24;
      opCodes[1001] <= 24;
      opCodes[1039] <= 24;
      opCodes[1077] <= 24;
      opCodes[1115] <= 24;
      opCodes[1155] <= 24;
      opCodes[1168] <= 24;
      opCodes[1199] <= 24;
      opCodes[1240] <= 24;
      opCodes[1251] <= 24;
      opCodes[1276] <= 24;
      opCodes[1314] <= 24;
      opCodes[1357] <= 24;
      opCodes[1370] <= 24;
      opCodes[1429] <= 24;
      opCodes[1440] <= 24;
      opCodes[1494] <= 24;
      opCodes[1532] <= 24;
      opCodes[1570] <= 24;
      opCodes[1608] <= 24;
      opCodes[1646] <= 24;
      opCodes[1659] <= 24;
      opCodes[1674] <= 24;
      opCodes[1727] <= 24;
      opCodes[1768] <= 24;
      opCodes[1779] <= 24;
      opCodes[1804] <= 24;
      opCodes[1842] <= 24;
      opCodes[1885] <= 24;
      opCodes[1898] <= 24;
      opCodes[1955] <= 24;
      opCodes[1966] <= 24;
      opCodes[2010] <= 24;
      opCodes[2051] <= 24;
      opCodes[2092] <= 24;
      opCodes[2133] <= 24;
      opCodes[2174] <= 24;
      opCodes[2215] <= 24;
      opCodes[2256] <= 24;
      opCodes[2297] <= 24;
      opCodes[2338] <= 24;
      opCodes[2379] <= 24;
      opCodes[2420] <= 24;
      opCodes[2461] <= 24;
      opCodes[2502] <= 24;
      opCodes[2543] <= 24;
      opCodes[2584] <= 24;
      opCodes[2625] <= 24;
      opCodes[2752] <= 24;
      opCodes[2765] <= 24;
      opCodes[2806] <= 24;
      opCodes[2847] <= 24;
      opCodes[2888] <= 24;
      opCodes[2929] <= 24;
      opCodes[2970] <= 24;
      opCodes[3011] <= 24;
      opCodes[3052] <= 24;
      opCodes[3093] <= 24;
      opCodes[3135] <= 24;
      opCodes[3158] <= 24;
      opCodes[3199] <= 24;
      opCodes[3240] <= 24;
      opCodes[3281] <= 24;
      opCodes[3322] <= 24;
      opCodes[3363] <= 24;
      opCodes[3404] <= 24;
      opCodes[3445] <= 24;
      opCodes[3486] <= 24;
      opCodes[3528] <= 24;
      opCodes[3651] <= 24;
      opCodes[3659] <= 24;
      opCodes[3706] <= 24;
      opCodes[3747] <= 24;
      opCodes[3788] <= 24;
      opCodes[3829] <= 24;
      opCodes[3870] <= 24;
      opCodes[3911] <= 24;
      opCodes[3952] <= 24;
      opCodes[3993] <= 24;
      opCodes[4061] <= 24;
      opCodes[4074] <= 24;
      opCodes[4114] <= 24;
      opCodes[4140] <= 24;
      opCodes[4181] <= 24;
      opCodes[4222] <= 24;
      opCodes[4263] <= 24;
      opCodes[4304] <= 24;
      opCodes[4345] <= 24;
      opCodes[4386] <= 24;
      opCodes[4427] <= 24;
      opCodes[4468] <= 24;
      opCodes[4543] <= 24;
      opCodes[4585] <= 24;
      opCodes[4596] <= 24;
      opCodes[4639] <= 24;
      opCodes[4680] <= 24;
      opCodes[4721] <= 24;
      opCodes[4762] <= 24;
      opCodes[4803] <= 24;
      opCodes[4844] <= 24;
      opCodes[4885] <= 24;
      opCodes[4926] <= 24;
      opCodes[4998] <= 24;
      opCodes[5008] <= 24;
      opCodes[5012] <= 24;
      opCodes[5038] <= 24;
      opCodes[5079] <= 24;
      opCodes[5120] <= 24;
      opCodes[5161] <= 24;
      opCodes[5202] <= 24;
      opCodes[5243] <= 24;
      opCodes[5284] <= 24;
      opCodes[5325] <= 24;
      opCodes[5366] <= 24;
      opCodes[5436] <= 24;
      opCodes[5444] <= 24;
      opCodes[5475] <= 24;
      opCodes[5516] <= 24;
      opCodes[5527] <= 24;
      opCodes[5599] <= 24;
      opCodes[5637] <= 24;
      opCodes[5675] <= 24;
      opCodes[5713] <= 24;
      opCodes[5751] <= 24;
      opCodes[5792] <= 24;
      opCodes[5843] <= 24;
      opCodes[5854] <= 24;
      opCodes[26] <= 25;
      opCodes[27] <= 26;
      opCodes[37] <= 26;
      opCodes[68] <= 26;
      opCodes[104] <= 26;
      opCodes[116] <= 26;
      opCodes[185] <= 26;
      opCodes[197] <= 26;
      opCodes[649] <= 26;
      opCodes[1201] <= 26;
      opCodes[1211] <= 26;
      opCodes[1242] <= 26;
      opCodes[1278] <= 26;
      opCodes[1290] <= 26;
      opCodes[1359] <= 26;
      opCodes[1371] <= 26;
      opCodes[1431] <= 26;
      opCodes[1453] <= 26;
      opCodes[1653] <= 26;
      opCodes[1677] <= 26;
      opCodes[1729] <= 26;
      opCodes[1739] <= 26;
      opCodes[1770] <= 26;
      opCodes[1806] <= 26;
      opCodes[1818] <= 26;
      opCodes[1887] <= 26;
      opCodes[1899] <= 26;
      opCodes[1960] <= 26;
      opCodes[3129] <= 26;
      opCodes[3522] <= 26;
      opCodes[3645] <= 26;
      opCodes[4055] <= 26;
      opCodes[4068] <= 26;
      opCodes[4528] <= 26;
      opCodes[4533] <= 26;
      opCodes[4590] <= 26;
      opCodes[4992] <= 26;
      opCodes[5430] <= 26;
      opCodes[5460] <= 26;
      opCodes[5465] <= 26;
      opCodes[5518] <= 26;
      opCodes[5558] <= 26;
      opCodes[5795] <= 26;
      opCodes[5845] <= 26;
      opCodes[28] <= 27;
      opCodes[69] <= 27;
      opCodes[105] <= 27;
      opCodes[126] <= 27;
      opCodes[150] <= 27;
      opCodes[186] <= 27;
      opCodes[224] <= 27;
      opCodes[352] <= 27;
      opCodes[355] <= 27;
      opCodes[370] <= 27;
      opCodes[390] <= 27;
      opCodes[393] <= 27;
      opCodes[408] <= 27;
      opCodes[428] <= 27;
      opCodes[431] <= 27;
      opCodes[446] <= 27;
      opCodes[466] <= 27;
      opCodes[469] <= 27;
      opCodes[484] <= 27;
      opCodes[504] <= 27;
      opCodes[507] <= 27;
      opCodes[522] <= 27;
      opCodes[542] <= 27;
      opCodes[545] <= 27;
      opCodes[560] <= 27;
      opCodes[580] <= 27;
      opCodes[583] <= 27;
      opCodes[598] <= 27;
      opCodes[618] <= 27;
      opCodes[621] <= 27;
      opCodes[636] <= 27;
      opCodes[680] <= 27;
      opCodes[693] <= 27;
      opCodes[781] <= 27;
      opCodes[784] <= 27;
      opCodes[799] <= 27;
      opCodes[819] <= 27;
      opCodes[822] <= 27;
      opCodes[837] <= 27;
      opCodes[857] <= 27;
      opCodes[860] <= 27;
      opCodes[875] <= 27;
      opCodes[895] <= 27;
      opCodes[898] <= 27;
      opCodes[913] <= 27;
      opCodes[933] <= 27;
      opCodes[936] <= 27;
      opCodes[955] <= 27;
      opCodes[975] <= 27;
      opCodes[978] <= 27;
      opCodes[993] <= 27;
      opCodes[1013] <= 27;
      opCodes[1016] <= 27;
      opCodes[1031] <= 27;
      opCodes[1051] <= 27;
      opCodes[1054] <= 27;
      opCodes[1069] <= 27;
      opCodes[1089] <= 27;
      opCodes[1092] <= 27;
      opCodes[1107] <= 27;
      opCodes[1127] <= 27;
      opCodes[1130] <= 27;
      opCodes[1147] <= 27;
      opCodes[1163] <= 27;
      opCodes[1176] <= 27;
      opCodes[1202] <= 27;
      opCodes[1243] <= 27;
      opCodes[1279] <= 27;
      opCodes[1300] <= 27;
      opCodes[1324] <= 27;
      opCodes[1360] <= 27;
      opCodes[1398] <= 27;
      opCodes[1432] <= 27;
      opCodes[1506] <= 27;
      opCodes[1509] <= 27;
      opCodes[1524] <= 27;
      opCodes[1544] <= 27;
      opCodes[1547] <= 27;
      opCodes[1562] <= 27;
      opCodes[1582] <= 27;
      opCodes[1585] <= 27;
      opCodes[1600] <= 27;
      opCodes[1620] <= 27;
      opCodes[1623] <= 27;
      opCodes[1638] <= 27;
      opCodes[1704] <= 27;
      opCodes[1730] <= 27;
      opCodes[1771] <= 27;
      opCodes[1807] <= 27;
      opCodes[1828] <= 27;
      opCodes[1852] <= 27;
      opCodes[1888] <= 27;
      opCodes[1926] <= 27;
      opCodes[2022] <= 27;
      opCodes[2025] <= 27;
      opCodes[2040] <= 27;
      opCodes[2063] <= 27;
      opCodes[2066] <= 27;
      opCodes[2081] <= 27;
      opCodes[2104] <= 27;
      opCodes[2107] <= 27;
      opCodes[2122] <= 27;
      opCodes[2145] <= 27;
      opCodes[2148] <= 27;
      opCodes[2163] <= 27;
      opCodes[2186] <= 27;
      opCodes[2189] <= 27;
      opCodes[2204] <= 27;
      opCodes[2227] <= 27;
      opCodes[2230] <= 27;
      opCodes[2245] <= 27;
      opCodes[2268] <= 27;
      opCodes[2271] <= 27;
      opCodes[2286] <= 27;
      opCodes[2309] <= 27;
      opCodes[2312] <= 27;
      opCodes[2327] <= 27;
      opCodes[2350] <= 27;
      opCodes[2353] <= 27;
      opCodes[2368] <= 27;
      opCodes[2391] <= 27;
      opCodes[2394] <= 27;
      opCodes[2409] <= 27;
      opCodes[2432] <= 27;
      opCodes[2435] <= 27;
      opCodes[2450] <= 27;
      opCodes[2473] <= 27;
      opCodes[2476] <= 27;
      opCodes[2491] <= 27;
      opCodes[2514] <= 27;
      opCodes[2517] <= 27;
      opCodes[2532] <= 27;
      opCodes[2555] <= 27;
      opCodes[2558] <= 27;
      opCodes[2573] <= 27;
      opCodes[2596] <= 27;
      opCodes[2599] <= 27;
      opCodes[2614] <= 27;
      opCodes[2637] <= 27;
      opCodes[2640] <= 27;
      opCodes[2655] <= 27;
      opCodes[2741] <= 27;
      opCodes[2777] <= 27;
      opCodes[2780] <= 27;
      opCodes[2795] <= 27;
      opCodes[2818] <= 27;
      opCodes[2821] <= 27;
      opCodes[2836] <= 27;
      opCodes[2859] <= 27;
      opCodes[2862] <= 27;
      opCodes[2877] <= 27;
      opCodes[2900] <= 27;
      opCodes[2903] <= 27;
      opCodes[2918] <= 27;
      opCodes[2941] <= 27;
      opCodes[2944] <= 27;
      opCodes[2959] <= 27;
      opCodes[2982] <= 27;
      opCodes[2985] <= 27;
      opCodes[3000] <= 27;
      opCodes[3023] <= 27;
      opCodes[3026] <= 27;
      opCodes[3041] <= 27;
      opCodes[3064] <= 27;
      opCodes[3067] <= 27;
      opCodes[3082] <= 27;
      opCodes[3105] <= 27;
      opCodes[3108] <= 27;
      opCodes[3123] <= 27;
      opCodes[3147] <= 27;
      opCodes[3170] <= 27;
      opCodes[3173] <= 27;
      opCodes[3188] <= 27;
      opCodes[3211] <= 27;
      opCodes[3214] <= 27;
      opCodes[3229] <= 27;
      opCodes[3252] <= 27;
      opCodes[3255] <= 27;
      opCodes[3270] <= 27;
      opCodes[3293] <= 27;
      opCodes[3296] <= 27;
      opCodes[3311] <= 27;
      opCodes[3334] <= 27;
      opCodes[3337] <= 27;
      opCodes[3352] <= 27;
      opCodes[3375] <= 27;
      opCodes[3378] <= 27;
      opCodes[3393] <= 27;
      opCodes[3416] <= 27;
      opCodes[3419] <= 27;
      opCodes[3434] <= 27;
      opCodes[3457] <= 27;
      opCodes[3460] <= 27;
      opCodes[3475] <= 27;
      opCodes[3498] <= 27;
      opCodes[3501] <= 27;
      opCodes[3516] <= 27;
      opCodes[3540] <= 27;
      opCodes[3618] <= 27;
      opCodes[3732] <= 27;
      opCodes[3773] <= 27;
      opCodes[3814] <= 27;
      opCodes[3855] <= 27;
      opCodes[3896] <= 27;
      opCodes[3937] <= 27;
      opCodes[3978] <= 27;
      opCodes[4019] <= 27;
      opCodes[4044] <= 27;
      opCodes[4102] <= 27;
      opCodes[4125] <= 27;
      opCodes[4166] <= 27;
      opCodes[4207] <= 27;
      opCodes[4248] <= 27;
      opCodes[4289] <= 27;
      opCodes[4330] <= 27;
      opCodes[4371] <= 27;
      opCodes[4412] <= 27;
      opCodes[4453] <= 27;
      opCodes[4494] <= 27;
      opCodes[4538] <= 27;
      opCodes[4551] <= 27;
      opCodes[4554] <= 27;
      opCodes[4591] <= 27;
      opCodes[4651] <= 27;
      opCodes[4654] <= 27;
      opCodes[4669] <= 27;
      opCodes[4692] <= 27;
      opCodes[4695] <= 27;
      opCodes[4710] <= 27;
      opCodes[4733] <= 27;
      opCodes[4736] <= 27;
      opCodes[4751] <= 27;
      opCodes[4774] <= 27;
      opCodes[4777] <= 27;
      opCodes[4792] <= 27;
      opCodes[4815] <= 27;
      opCodes[4818] <= 27;
      opCodes[4833] <= 27;
      opCodes[4856] <= 27;
      opCodes[4859] <= 27;
      opCodes[4874] <= 27;
      opCodes[4897] <= 27;
      opCodes[4900] <= 27;
      opCodes[4915] <= 27;
      opCodes[4938] <= 27;
      opCodes[4941] <= 27;
      opCodes[4956] <= 27;
      opCodes[4981] <= 27;
      opCodes[5022] <= 27;
      opCodes[5027] <= 27;
      opCodes[5050] <= 27;
      opCodes[5053] <= 27;
      opCodes[5068] <= 27;
      opCodes[5091] <= 27;
      opCodes[5094] <= 27;
      opCodes[5109] <= 27;
      opCodes[5132] <= 27;
      opCodes[5135] <= 27;
      opCodes[5150] <= 27;
      opCodes[5173] <= 27;
      opCodes[5176] <= 27;
      opCodes[5191] <= 27;
      opCodes[5214] <= 27;
      opCodes[5217] <= 27;
      opCodes[5232] <= 27;
      opCodes[5255] <= 27;
      opCodes[5258] <= 27;
      opCodes[5273] <= 27;
      opCodes[5296] <= 27;
      opCodes[5299] <= 27;
      opCodes[5314] <= 27;
      opCodes[5337] <= 27;
      opCodes[5340] <= 27;
      opCodes[5355] <= 27;
      opCodes[5378] <= 27;
      opCodes[5381] <= 27;
      opCodes[5396] <= 27;
      opCodes[5431] <= 27;
      opCodes[5456] <= 27;
      opCodes[5461] <= 27;
      opCodes[5470] <= 27;
      opCodes[5483] <= 27;
      opCodes[5486] <= 27;
      opCodes[5494] <= 27;
      opCodes[5519] <= 27;
      opCodes[5531] <= 27;
      opCodes[5611] <= 27;
      opCodes[5614] <= 27;
      opCodes[5629] <= 27;
      opCodes[5649] <= 27;
      opCodes[5652] <= 27;
      opCodes[5667] <= 27;
      opCodes[5687] <= 27;
      opCodes[5690] <= 27;
      opCodes[5705] <= 27;
      opCodes[5725] <= 27;
      opCodes[5728] <= 27;
      opCodes[5743] <= 27;
      opCodes[5763] <= 27;
      opCodes[5766] <= 27;
      opCodes[5785] <= 27;
      opCodes[5822] <= 27;
      opCodes[5846] <= 27;
      opCodes[5862] <= 27;
      opCodes[29] <= 28;
      opCodes[70] <= 28;
      opCodes[106] <= 28;
      opCodes[142] <= 28;
      opCodes[187] <= 28;
      opCodes[364] <= 28;
      opCodes[402] <= 28;
      opCodes[440] <= 28;
      opCodes[478] <= 28;
      opCodes[516] <= 28;
      opCodes[554] <= 28;
      opCodes[592] <= 28;
      opCodes[630] <= 28;
      opCodes[648] <= 28;
      opCodes[651] <= 28;
      opCodes[674] <= 28;
      opCodes[687] <= 28;
      opCodes[793] <= 28;
      opCodes[831] <= 28;
      opCodes[869] <= 28;
      opCodes[907] <= 28;
      opCodes[949] <= 28;
      opCodes[987] <= 28;
      opCodes[1025] <= 28;
      opCodes[1063] <= 28;
      opCodes[1101] <= 28;
      opCodes[1141] <= 28;
      opCodes[1157] <= 28;
      opCodes[1170] <= 28;
      opCodes[1203] <= 28;
      opCodes[1244] <= 28;
      opCodes[1280] <= 28;
      opCodes[1316] <= 28;
      opCodes[1361] <= 28;
      opCodes[1433] <= 28;
      opCodes[1518] <= 28;
      opCodes[1556] <= 28;
      opCodes[1594] <= 28;
      opCodes[1632] <= 28;
      opCodes[1652] <= 28;
      opCodes[1655] <= 28;
      opCodes[1676] <= 28;
      opCodes[1731] <= 28;
      opCodes[1772] <= 28;
      opCodes[1808] <= 28;
      opCodes[1844] <= 28;
      opCodes[1889] <= 28;
      opCodes[1959] <= 28;
      opCodes[1962] <= 28;
      opCodes[2034] <= 28;
      opCodes[2075] <= 28;
      opCodes[2116] <= 28;
      opCodes[2157] <= 28;
      opCodes[2198] <= 28;
      opCodes[2239] <= 28;
      opCodes[2280] <= 28;
      opCodes[2321] <= 28;
      opCodes[2362] <= 28;
      opCodes[2403] <= 28;
      opCodes[2444] <= 28;
      opCodes[2485] <= 28;
      opCodes[2526] <= 28;
      opCodes[2567] <= 28;
      opCodes[2608] <= 28;
      opCodes[2649] <= 28;
      opCodes[2789] <= 28;
      opCodes[2830] <= 28;
      opCodes[2871] <= 28;
      opCodes[2912] <= 28;
      opCodes[2953] <= 28;
      opCodes[2994] <= 28;
      opCodes[3035] <= 28;
      opCodes[3076] <= 28;
      opCodes[3117] <= 28;
      opCodes[3128] <= 28;
      opCodes[3131] <= 28;
      opCodes[3141] <= 28;
      opCodes[3182] <= 28;
      opCodes[3223] <= 28;
      opCodes[3264] <= 28;
      opCodes[3305] <= 28;
      opCodes[3346] <= 28;
      opCodes[3387] <= 28;
      opCodes[3428] <= 28;
      opCodes[3469] <= 28;
      opCodes[3510] <= 28;
      opCodes[3521] <= 28;
      opCodes[3524] <= 28;
      opCodes[3534] <= 28;
      opCodes[3644] <= 28;
      opCodes[3647] <= 28;
      opCodes[3655] <= 28;
      opCodes[3702] <= 28;
      opCodes[3743] <= 28;
      opCodes[3784] <= 28;
      opCodes[3825] <= 28;
      opCodes[3866] <= 28;
      opCodes[3907] <= 28;
      opCodes[3948] <= 28;
      opCodes[3989] <= 28;
      opCodes[4054] <= 28;
      opCodes[4057] <= 28;
      opCodes[4067] <= 28;
      opCodes[4070] <= 28;
      opCodes[4110] <= 28;
      opCodes[4136] <= 28;
      opCodes[4177] <= 28;
      opCodes[4218] <= 28;
      opCodes[4259] <= 28;
      opCodes[4300] <= 28;
      opCodes[4341] <= 28;
      opCodes[4382] <= 28;
      opCodes[4423] <= 28;
      opCodes[4464] <= 28;
      opCodes[4527] <= 28;
      opCodes[4530] <= 28;
      opCodes[4581] <= 28;
      opCodes[4589] <= 28;
      opCodes[4592] <= 28;
      opCodes[4663] <= 28;
      opCodes[4704] <= 28;
      opCodes[4745] <= 28;
      opCodes[4786] <= 28;
      opCodes[4827] <= 28;
      opCodes[4868] <= 28;
      opCodes[4909] <= 28;
      opCodes[4950] <= 28;
      opCodes[4991] <= 28;
      opCodes[4994] <= 28;
      opCodes[5004] <= 28;
      opCodes[5014] <= 28;
      opCodes[5062] <= 28;
      opCodes[5103] <= 28;
      opCodes[5144] <= 28;
      opCodes[5185] <= 28;
      opCodes[5226] <= 28;
      opCodes[5267] <= 28;
      opCodes[5308] <= 28;
      opCodes[5349] <= 28;
      opCodes[5390] <= 28;
      opCodes[5429] <= 28;
      opCodes[5432] <= 28;
      opCodes[5440] <= 28;
      opCodes[5448] <= 28;
      opCodes[5459] <= 28;
      opCodes[5462] <= 28;
      opCodes[5520] <= 28;
      opCodes[5623] <= 28;
      opCodes[5661] <= 28;
      opCodes[5699] <= 28;
      opCodes[5737] <= 28;
      opCodes[5779] <= 28;
      opCodes[5794] <= 28;
      opCodes[5847] <= 28;
      opCodes[32] <= 29;
      opCodes[33] <= 30;
      opCodes[44] <= 30;
      opCodes[334] <= 30;
      opCodes[372] <= 30;
      opCodes[410] <= 30;
      opCodes[448] <= 30;
      opCodes[486] <= 30;
      opCodes[524] <= 30;
      opCodes[562] <= 30;
      opCodes[600] <= 30;
      opCodes[666] <= 30;
      opCodes[682] <= 30;
      opCodes[763] <= 30;
      opCodes[801] <= 30;
      opCodes[839] <= 30;
      opCodes[877] <= 30;
      opCodes[915] <= 30;
      opCodes[946] <= 30;
      opCodes[957] <= 30;
      opCodes[995] <= 30;
      opCodes[1033] <= 30;
      opCodes[1071] <= 30;
      opCodes[1109] <= 30;
      opCodes[1138] <= 30;
      opCodes[1149] <= 30;
      opCodes[1165] <= 30;
      opCodes[1207] <= 30;
      opCodes[1218] <= 30;
      opCodes[1407] <= 30;
      opCodes[1735] <= 30;
      opCodes[1746] <= 30;
      opCodes[1969] <= 30;
      opCodes[1998] <= 30;
      opCodes[2031] <= 30;
      opCodes[2072] <= 30;
      opCodes[2113] <= 30;
      opCodes[2154] <= 30;
      opCodes[2195] <= 30;
      opCodes[2236] <= 30;
      opCodes[2277] <= 30;
      opCodes[2318] <= 30;
      opCodes[2359] <= 30;
      opCodes[2400] <= 30;
      opCodes[2441] <= 30;
      opCodes[2482] <= 30;
      opCodes[2523] <= 30;
      opCodes[2564] <= 30;
      opCodes[2605] <= 30;
      opCodes[2646] <= 30;
      opCodes[2657] <= 30;
      opCodes[2746] <= 30;
      opCodes[2786] <= 30;
      opCodes[2827] <= 30;
      opCodes[2868] <= 30;
      opCodes[2909] <= 30;
      opCodes[2950] <= 30;
      opCodes[2991] <= 30;
      opCodes[3032] <= 30;
      opCodes[3073] <= 30;
      opCodes[3114] <= 30;
      opCodes[3136] <= 30;
      opCodes[3179] <= 30;
      opCodes[3220] <= 30;
      opCodes[3261] <= 30;
      opCodes[3302] <= 30;
      opCodes[3343] <= 30;
      opCodes[3384] <= 30;
      opCodes[3425] <= 30;
      opCodes[3466] <= 30;
      opCodes[3507] <= 30;
      opCodes[3529] <= 30;
      opCodes[3531] <= 30;
      opCodes[3598] <= 30;
      opCodes[5776] <= 30;
      opCodes[34] <= 31;
      opCodes[113] <= 31;
      opCodes[1208] <= 31;
      opCodes[1287] <= 31;
      opCodes[1736] <= 31;
      opCodes[1815] <= 31;
      opCodes[35] <= 32;
      opCodes[114] <= 32;
      opCodes[1209] <= 32;
      opCodes[1288] <= 32;
      opCodes[1737] <= 32;
      opCodes[1816] <= 32;
      opCodes[36] <= 33;
      opCodes[115] <= 33;
      opCodes[1210] <= 33;
      opCodes[1289] <= 33;
      opCodes[1738] <= 33;
      opCodes[1817] <= 33;
      opCodes[38] <= 34;
      opCodes[117] <= 34;
      opCodes[1212] <= 34;
      opCodes[1291] <= 34;
      opCodes[1740] <= 34;
      opCodes[1819] <= 34;
      opCodes[39] <= 35;
      opCodes[118] <= 35;
      opCodes[143] <= 35;
      opCodes[219] <= 35;
      opCodes[365] <= 35;
      opCodes[403] <= 35;
      opCodes[441] <= 35;
      opCodes[479] <= 35;
      opCodes[517] <= 35;
      opCodes[555] <= 35;
      opCodes[593] <= 35;
      opCodes[631] <= 35;
      opCodes[643] <= 35;
      opCodes[656] <= 35;
      opCodes[675] <= 35;
      opCodes[688] <= 35;
      opCodes[794] <= 35;
      opCodes[832] <= 35;
      opCodes[870] <= 35;
      opCodes[908] <= 35;
      opCodes[942] <= 35;
      opCodes[950] <= 35;
      opCodes[988] <= 35;
      opCodes[1026] <= 35;
      opCodes[1064] <= 35;
      opCodes[1102] <= 35;
      opCodes[1142] <= 35;
      opCodes[1158] <= 35;
      opCodes[1171] <= 35;
      opCodes[1213] <= 35;
      opCodes[1292] <= 35;
      opCodes[1317] <= 35;
      opCodes[1393] <= 35;
      opCodes[1519] <= 35;
      opCodes[1557] <= 35;
      opCodes[1595] <= 35;
      opCodes[1633] <= 35;
      opCodes[1647] <= 35;
      opCodes[1660] <= 35;
      opCodes[1699] <= 35;
      opCodes[1741] <= 35;
      opCodes[1820] <= 35;
      opCodes[1845] <= 35;
      opCodes[1921] <= 35;
      opCodes[2035] <= 35;
      opCodes[2076] <= 35;
      opCodes[2117] <= 35;
      opCodes[2158] <= 35;
      opCodes[2199] <= 35;
      opCodes[2240] <= 35;
      opCodes[2281] <= 35;
      opCodes[2322] <= 35;
      opCodes[2363] <= 35;
      opCodes[2404] <= 35;
      opCodes[2445] <= 35;
      opCodes[2486] <= 35;
      opCodes[2527] <= 35;
      opCodes[2568] <= 35;
      opCodes[2609] <= 35;
      opCodes[2650] <= 35;
      opCodes[2753] <= 35;
      opCodes[2790] <= 35;
      opCodes[2831] <= 35;
      opCodes[2872] <= 35;
      opCodes[2913] <= 35;
      opCodes[2954] <= 35;
      opCodes[2995] <= 35;
      opCodes[3036] <= 35;
      opCodes[3077] <= 35;
      opCodes[3118] <= 35;
      opCodes[3142] <= 35;
      opCodes[3183] <= 35;
      opCodes[3224] <= 35;
      opCodes[3265] <= 35;
      opCodes[3306] <= 35;
      opCodes[3347] <= 35;
      opCodes[3388] <= 35;
      opCodes[3429] <= 35;
      opCodes[3470] <= 35;
      opCodes[3511] <= 35;
      opCodes[3535] <= 35;
      opCodes[3727] <= 35;
      opCodes[3768] <= 35;
      opCodes[3809] <= 35;
      opCodes[3850] <= 35;
      opCodes[3891] <= 35;
      opCodes[3932] <= 35;
      opCodes[3973] <= 35;
      opCodes[4014] <= 35;
      opCodes[4062] <= 35;
      opCodes[4097] <= 35;
      opCodes[4161] <= 35;
      opCodes[4202] <= 35;
      opCodes[4243] <= 35;
      opCodes[4284] <= 35;
      opCodes[4325] <= 35;
      opCodes[4366] <= 35;
      opCodes[4407] <= 35;
      opCodes[4448] <= 35;
      opCodes[4489] <= 35;
      opCodes[4664] <= 35;
      opCodes[4705] <= 35;
      opCodes[4746] <= 35;
      opCodes[4787] <= 35;
      opCodes[4828] <= 35;
      opCodes[4869] <= 35;
      opCodes[4910] <= 35;
      opCodes[4951] <= 35;
      opCodes[5015] <= 35;
      opCodes[5063] <= 35;
      opCodes[5104] <= 35;
      opCodes[5145] <= 35;
      opCodes[5186] <= 35;
      opCodes[5227] <= 35;
      opCodes[5268] <= 35;
      opCodes[5309] <= 35;
      opCodes[5350] <= 35;
      opCodes[5391] <= 35;
      opCodes[5437] <= 35;
      opCodes[5449] <= 35;
      opCodes[5624] <= 35;
      opCodes[5662] <= 35;
      opCodes[5700] <= 35;
      opCodes[5738] <= 35;
      opCodes[5772] <= 35;
      opCodes[5780] <= 35;
      opCodes[5817] <= 35;
      opCodes[40] <= 36;
      opCodes[119] <= 36;
      opCodes[1214] <= 36;
      opCodes[1293] <= 36;
      opCodes[1742] <= 36;
      opCodes[1821] <= 36;
      opCodes[41] <= 37;
      opCodes[78] <= 37;
      opCodes[120] <= 37;
      opCodes[145] <= 37;
      opCodes[221] <= 37;
      opCodes[367] <= 37;
      opCodes[405] <= 37;
      opCodes[443] <= 37;
      opCodes[481] <= 37;
      opCodes[519] <= 37;
      opCodes[557] <= 37;
      opCodes[595] <= 37;
      opCodes[633] <= 37;
      opCodes[677] <= 37;
      opCodes[690] <= 37;
      opCodes[796] <= 37;
      opCodes[834] <= 37;
      opCodes[872] <= 37;
      opCodes[910] <= 37;
      opCodes[952] <= 37;
      opCodes[990] <= 37;
      opCodes[1028] <= 37;
      opCodes[1066] <= 37;
      opCodes[1104] <= 37;
      opCodes[1144] <= 37;
      opCodes[1160] <= 37;
      opCodes[1173] <= 37;
      opCodes[1215] <= 37;
      opCodes[1252] <= 37;
      opCodes[1294] <= 37;
      opCodes[1319] <= 37;
      opCodes[1395] <= 37;
      opCodes[1441] <= 37;
      opCodes[1521] <= 37;
      opCodes[1559] <= 37;
      opCodes[1597] <= 37;
      opCodes[1635] <= 37;
      opCodes[1701] <= 37;
      opCodes[1743] <= 37;
      opCodes[1780] <= 37;
      opCodes[1822] <= 37;
      opCodes[1847] <= 37;
      opCodes[1923] <= 37;
      opCodes[1956] <= 37;
      opCodes[1967] <= 37;
      opCodes[2037] <= 37;
      opCodes[2078] <= 37;
      opCodes[2119] <= 37;
      opCodes[2160] <= 37;
      opCodes[2201] <= 37;
      opCodes[2242] <= 37;
      opCodes[2283] <= 37;
      opCodes[2324] <= 37;
      opCodes[2365] <= 37;
      opCodes[2406] <= 37;
      opCodes[2447] <= 37;
      opCodes[2488] <= 37;
      opCodes[2529] <= 37;
      opCodes[2570] <= 37;
      opCodes[2611] <= 37;
      opCodes[2652] <= 37;
      opCodes[2792] <= 37;
      opCodes[2833] <= 37;
      opCodes[2874] <= 37;
      opCodes[2915] <= 37;
      opCodes[2956] <= 37;
      opCodes[2997] <= 37;
      opCodes[3038] <= 37;
      opCodes[3079] <= 37;
      opCodes[3120] <= 37;
      opCodes[3144] <= 37;
      opCodes[3185] <= 37;
      opCodes[3226] <= 37;
      opCodes[3267] <= 37;
      opCodes[3308] <= 37;
      opCodes[3349] <= 37;
      opCodes[3390] <= 37;
      opCodes[3431] <= 37;
      opCodes[3472] <= 37;
      opCodes[3513] <= 37;
      opCodes[3537] <= 37;
      opCodes[3652] <= 37;
      opCodes[3660] <= 37;
      opCodes[3729] <= 37;
      opCodes[3770] <= 37;
      opCodes[3811] <= 37;
      opCodes[3852] <= 37;
      opCodes[3893] <= 37;
      opCodes[3934] <= 37;
      opCodes[3975] <= 37;
      opCodes[4016] <= 37;
      opCodes[4099] <= 37;
      opCodes[4163] <= 37;
      opCodes[4204] <= 37;
      opCodes[4245] <= 37;
      opCodes[4286] <= 37;
      opCodes[4327] <= 37;
      opCodes[4368] <= 37;
      opCodes[4409] <= 37;
      opCodes[4450] <= 37;
      opCodes[4491] <= 37;
      opCodes[4586] <= 37;
      opCodes[4597] <= 37;
      opCodes[4666] <= 37;
      opCodes[4707] <= 37;
      opCodes[4748] <= 37;
      opCodes[4789] <= 37;
      opCodes[4830] <= 37;
      opCodes[4871] <= 37;
      opCodes[4912] <= 37;
      opCodes[4953] <= 37;
      opCodes[4999] <= 37;
      opCodes[5017] <= 37;
      opCodes[5065] <= 37;
      opCodes[5106] <= 37;
      opCodes[5147] <= 37;
      opCodes[5188] <= 37;
      opCodes[5229] <= 37;
      opCodes[5270] <= 37;
      opCodes[5311] <= 37;
      opCodes[5352] <= 37;
      opCodes[5393] <= 37;
      opCodes[5451] <= 37;
      opCodes[5528] <= 37;
      opCodes[5626] <= 37;
      opCodes[5664] <= 37;
      opCodes[5702] <= 37;
      opCodes[5740] <= 37;
      opCodes[5782] <= 37;
      opCodes[5819] <= 37;
      opCodes[5855] <= 37;
      opCodes[42] <= 38;
      opCodes[121] <= 38;
      opCodes[1216] <= 38;
      opCodes[1295] <= 38;
      opCodes[1744] <= 38;
      opCodes[1823] <= 38;
      opCodes[43] <= 39;
      opCodes[122] <= 39;
      opCodes[45] <= 40;
      opCodes[124] <= 40;
      opCodes[1219] <= 40;
      opCodes[1298] <= 40;
      opCodes[1408] <= 40;
      opCodes[1747] <= 40;
      opCodes[1826] <= 40;
      opCodes[3599] <= 40;
      opCodes[5529] <= 40;
      opCodes[5856] <= 40;
      opCodes[5860] <= 40;
      opCodes[46] <= 41;
      opCodes[1220] <= 41;
      opCodes[1748] <= 41;
      opCodes[47] <= 42;
      opCodes[1221] <= 42;
      opCodes[1410] <= 42;
      opCodes[1451] <= 42;
      opCodes[1749] <= 42;
      opCodes[3602] <= 42;
      opCodes[3608] <= 42;
      opCodes[3623] <= 42;
      opCodes[4566] <= 42;
      opCodes[5497] <= 42;
      opCodes[5556] <= 42;
      opCodes[5824] <= 42;
      opCodes[48] <= 43;
      opCodes[87] <= 43;
      opCodes[136] <= 43;
      opCodes[168] <= 43;
      opCodes[192] <= 43;
      opCodes[335] <= 43;
      opCodes[362] <= 43;
      opCodes[373] <= 43;
      opCodes[400] <= 43;
      opCodes[411] <= 43;
      opCodes[438] <= 43;
      opCodes[449] <= 43;
      opCodes[476] <= 43;
      opCodes[487] <= 43;
      opCodes[514] <= 43;
      opCodes[525] <= 43;
      opCodes[552] <= 43;
      opCodes[563] <= 43;
      opCodes[590] <= 43;
      opCodes[601] <= 43;
      opCodes[628] <= 43;
      opCodes[646] <= 43;
      opCodes[667] <= 43;
      opCodes[764] <= 43;
      opCodes[791] <= 43;
      opCodes[802] <= 43;
      opCodes[829] <= 43;
      opCodes[840] <= 43;
      opCodes[867] <= 43;
      opCodes[878] <= 43;
      opCodes[905] <= 43;
      opCodes[916] <= 43;
      opCodes[945] <= 43;
      opCodes[958] <= 43;
      opCodes[985] <= 43;
      opCodes[996] <= 43;
      opCodes[1023] <= 43;
      opCodes[1034] <= 43;
      opCodes[1061] <= 43;
      opCodes[1072] <= 43;
      opCodes[1099] <= 43;
      opCodes[1110] <= 43;
      opCodes[1137] <= 43;
      opCodes[1150] <= 43;
      opCodes[1222] <= 43;
      opCodes[1261] <= 43;
      opCodes[1310] <= 43;
      opCodes[1342] <= 43;
      opCodes[1366] <= 43;
      opCodes[1411] <= 43;
      opCodes[1489] <= 43;
      opCodes[1516] <= 43;
      opCodes[1527] <= 43;
      opCodes[1554] <= 43;
      opCodes[1565] <= 43;
      opCodes[1592] <= 43;
      opCodes[1603] <= 43;
      opCodes[1630] <= 43;
      opCodes[1641] <= 43;
      opCodes[1650] <= 43;
      opCodes[1670] <= 43;
      opCodes[1750] <= 43;
      opCodes[1789] <= 43;
      opCodes[1838] <= 43;
      opCodes[1870] <= 43;
      opCodes[1894] <= 43;
      opCodes[1999] <= 43;
      opCodes[2005] <= 43;
      opCodes[2032] <= 43;
      opCodes[2046] <= 43;
      opCodes[2073] <= 43;
      opCodes[2087] <= 43;
      opCodes[2114] <= 43;
      opCodes[2128] <= 43;
      opCodes[2155] <= 43;
      opCodes[2169] <= 43;
      opCodes[2196] <= 43;
      opCodes[2210] <= 43;
      opCodes[2237] <= 43;
      opCodes[2251] <= 43;
      opCodes[2278] <= 43;
      opCodes[2292] <= 43;
      opCodes[2319] <= 43;
      opCodes[2333] <= 43;
      opCodes[2360] <= 43;
      opCodes[2374] <= 43;
      opCodes[2401] <= 43;
      opCodes[2415] <= 43;
      opCodes[2442] <= 43;
      opCodes[2456] <= 43;
      opCodes[2483] <= 43;
      opCodes[2497] <= 43;
      opCodes[2524] <= 43;
      opCodes[2538] <= 43;
      opCodes[2565] <= 43;
      opCodes[2579] <= 43;
      opCodes[2606] <= 43;
      opCodes[2620] <= 43;
      opCodes[2647] <= 43;
      opCodes[2747] <= 43;
      opCodes[2760] <= 43;
      opCodes[2787] <= 43;
      opCodes[2801] <= 43;
      opCodes[2828] <= 43;
      opCodes[2842] <= 43;
      opCodes[2869] <= 43;
      opCodes[2883] <= 43;
      opCodes[2910] <= 43;
      opCodes[2924] <= 43;
      opCodes[2951] <= 43;
      opCodes[2965] <= 43;
      opCodes[2992] <= 43;
      opCodes[3006] <= 43;
      opCodes[3033] <= 43;
      opCodes[3047] <= 43;
      opCodes[3074] <= 43;
      opCodes[3088] <= 43;
      opCodes[3115] <= 43;
      opCodes[3126] <= 43;
      opCodes[3137] <= 43;
      opCodes[3153] <= 43;
      opCodes[3180] <= 43;
      opCodes[3194] <= 43;
      opCodes[3221] <= 43;
      opCodes[3235] <= 43;
      opCodes[3262] <= 43;
      opCodes[3276] <= 43;
      opCodes[3303] <= 43;
      opCodes[3317] <= 43;
      opCodes[3344] <= 43;
      opCodes[3358] <= 43;
      opCodes[3385] <= 43;
      opCodes[3399] <= 43;
      opCodes[3426] <= 43;
      opCodes[3440] <= 43;
      opCodes[3467] <= 43;
      opCodes[3481] <= 43;
      opCodes[3508] <= 43;
      opCodes[3519] <= 43;
      opCodes[3530] <= 43;
      opCodes[3642] <= 43;
      opCodes[3697] <= 43;
      opCodes[3708] <= 43;
      opCodes[3738] <= 43;
      opCodes[3749] <= 43;
      opCodes[3779] <= 43;
      opCodes[3790] <= 43;
      opCodes[3820] <= 43;
      opCodes[3831] <= 43;
      opCodes[3861] <= 43;
      opCodes[3872] <= 43;
      opCodes[3902] <= 43;
      opCodes[3913] <= 43;
      opCodes[3943] <= 43;
      opCodes[3954] <= 43;
      opCodes[3984] <= 43;
      opCodes[3995] <= 43;
      opCodes[4052] <= 43;
      opCodes[4065] <= 43;
      opCodes[4076] <= 43;
      opCodes[4105] <= 43;
      opCodes[4131] <= 43;
      opCodes[4142] <= 43;
      opCodes[4172] <= 43;
      opCodes[4183] <= 43;
      opCodes[4213] <= 43;
      opCodes[4224] <= 43;
      opCodes[4254] <= 43;
      opCodes[4265] <= 43;
      opCodes[4295] <= 43;
      opCodes[4306] <= 43;
      opCodes[4336] <= 43;
      opCodes[4347] <= 43;
      opCodes[4377] <= 43;
      opCodes[4388] <= 43;
      opCodes[4418] <= 43;
      opCodes[4429] <= 43;
      opCodes[4459] <= 43;
      opCodes[4470] <= 43;
      opCodes[4525] <= 43;
      opCodes[4579] <= 43;
      opCodes[4634] <= 43;
      opCodes[4661] <= 43;
      opCodes[4675] <= 43;
      opCodes[4702] <= 43;
      opCodes[4716] <= 43;
      opCodes[4743] <= 43;
      opCodes[4757] <= 43;
      opCodes[4784] <= 43;
      opCodes[4798] <= 43;
      opCodes[4825] <= 43;
      opCodes[4839] <= 43;
      opCodes[4866] <= 43;
      opCodes[4880] <= 43;
      opCodes[4907] <= 43;
      opCodes[4921] <= 43;
      opCodes[4948] <= 43;
      opCodes[4989] <= 43;
      opCodes[5002] <= 43;
      opCodes[5010] <= 43;
      opCodes[5033] <= 43;
      opCodes[5060] <= 43;
      opCodes[5074] <= 43;
      opCodes[5101] <= 43;
      opCodes[5115] <= 43;
      opCodes[5142] <= 43;
      opCodes[5156] <= 43;
      opCodes[5183] <= 43;
      opCodes[5197] <= 43;
      opCodes[5224] <= 43;
      opCodes[5238] <= 43;
      opCodes[5265] <= 43;
      opCodes[5279] <= 43;
      opCodes[5306] <= 43;
      opCodes[5320] <= 43;
      opCodes[5347] <= 43;
      opCodes[5361] <= 43;
      opCodes[5388] <= 43;
      opCodes[5427] <= 43;
      opCodes[5498] <= 43;
      opCodes[5594] <= 43;
      opCodes[5621] <= 43;
      opCodes[5632] <= 43;
      opCodes[5659] <= 43;
      opCodes[5670] <= 43;
      opCodes[5697] <= 43;
      opCodes[5708] <= 43;
      opCodes[5735] <= 43;
      opCodes[5746] <= 43;
      opCodes[5775] <= 43;
      opCodes[5788] <= 43;
      opCodes[5825] <= 43;
      opCodes[55] <= 44;
      opCodes[1229] <= 44;
      opCodes[1418] <= 44;
      opCodes[1757] <= 44;
      opCodes[5505] <= 44;
      opCodes[5832] <= 44;
      opCodes[56] <= 45;
      opCodes[204] <= 45;
      opCodes[213] <= 45;
      opCodes[216] <= 45;
      opCodes[254] <= 45;
      opCodes[359] <= 45;
      opCodes[397] <= 45;
      opCodes[435] <= 45;
      opCodes[473] <= 45;
      opCodes[511] <= 45;
      opCodes[549] <= 45;
      opCodes[587] <= 45;
      opCodes[625] <= 45;
      opCodes[650] <= 45;
      opCodes[788] <= 45;
      opCodes[826] <= 45;
      opCodes[864] <= 45;
      opCodes[902] <= 45;
      opCodes[940] <= 45;
      opCodes[982] <= 45;
      opCodes[1020] <= 45;
      opCodes[1058] <= 45;
      opCodes[1096] <= 45;
      opCodes[1134] <= 45;
      opCodes[1230] <= 45;
      opCodes[1378] <= 45;
      opCodes[1387] <= 45;
      opCodes[1390] <= 45;
      opCodes[1419] <= 45;
      opCodes[1513] <= 45;
      opCodes[1551] <= 45;
      opCodes[1589] <= 45;
      opCodes[1627] <= 45;
      opCodes[1654] <= 45;
      opCodes[1684] <= 45;
      opCodes[1693] <= 45;
      opCodes[1696] <= 45;
      opCodes[1758] <= 45;
      opCodes[1906] <= 45;
      opCodes[1915] <= 45;
      opCodes[1918] <= 45;
      opCodes[1943] <= 45;
      opCodes[1961] <= 45;
      opCodes[2029] <= 45;
      opCodes[2070] <= 45;
      opCodes[2111] <= 45;
      opCodes[2152] <= 45;
      opCodes[2193] <= 45;
      opCodes[2234] <= 45;
      opCodes[2275] <= 45;
      opCodes[2316] <= 45;
      opCodes[2357] <= 45;
      opCodes[2398] <= 45;
      opCodes[2439] <= 45;
      opCodes[2480] <= 45;
      opCodes[2521] <= 45;
      opCodes[2562] <= 45;
      opCodes[2603] <= 45;
      opCodes[2644] <= 45;
      opCodes[2723] <= 45;
      opCodes[2732] <= 45;
      opCodes[2784] <= 45;
      opCodes[2825] <= 45;
      opCodes[2866] <= 45;
      opCodes[2907] <= 45;
      opCodes[2948] <= 45;
      opCodes[2989] <= 45;
      opCodes[3030] <= 45;
      opCodes[3071] <= 45;
      opCodes[3112] <= 45;
      opCodes[3130] <= 45;
      opCodes[3177] <= 45;
      opCodes[3218] <= 45;
      opCodes[3259] <= 45;
      opCodes[3300] <= 45;
      opCodes[3341] <= 45;
      opCodes[3382] <= 45;
      opCodes[3423] <= 45;
      opCodes[3464] <= 45;
      opCodes[3505] <= 45;
      opCodes[3523] <= 45;
      opCodes[3613] <= 45;
      opCodes[3635] <= 45;
      opCodes[3646] <= 45;
      opCodes[3699] <= 45;
      opCodes[3716] <= 45;
      opCodes[3723] <= 45;
      opCodes[3740] <= 45;
      opCodes[3757] <= 45;
      opCodes[3764] <= 45;
      opCodes[3781] <= 45;
      opCodes[3798] <= 45;
      opCodes[3805] <= 45;
      opCodes[3822] <= 45;
      opCodes[3839] <= 45;
      opCodes[3846] <= 45;
      opCodes[3863] <= 45;
      opCodes[3880] <= 45;
      opCodes[3887] <= 45;
      opCodes[3904] <= 45;
      opCodes[3921] <= 45;
      opCodes[3928] <= 45;
      opCodes[3945] <= 45;
      opCodes[3962] <= 45;
      opCodes[3969] <= 45;
      opCodes[3986] <= 45;
      opCodes[4003] <= 45;
      opCodes[4010] <= 45;
      opCodes[4028] <= 45;
      opCodes[4037] <= 45;
      opCodes[4056] <= 45;
      opCodes[4069] <= 45;
      opCodes[4086] <= 45;
      opCodes[4093] <= 45;
      opCodes[4107] <= 45;
      opCodes[4120] <= 45;
      opCodes[4133] <= 45;
      opCodes[4150] <= 45;
      opCodes[4157] <= 45;
      opCodes[4174] <= 45;
      opCodes[4191] <= 45;
      opCodes[4198] <= 45;
      opCodes[4215] <= 45;
      opCodes[4232] <= 45;
      opCodes[4239] <= 45;
      opCodes[4256] <= 45;
      opCodes[4273] <= 45;
      opCodes[4280] <= 45;
      opCodes[4297] <= 45;
      opCodes[4314] <= 45;
      opCodes[4321] <= 45;
      opCodes[4338] <= 45;
      opCodes[4355] <= 45;
      opCodes[4362] <= 45;
      opCodes[4379] <= 45;
      opCodes[4396] <= 45;
      opCodes[4403] <= 45;
      opCodes[4420] <= 45;
      opCodes[4437] <= 45;
      opCodes[4444] <= 45;
      opCodes[4461] <= 45;
      opCodes[4478] <= 45;
      opCodes[4485] <= 45;
      opCodes[4529] <= 45;
      opCodes[4558] <= 45;
      opCodes[4564] <= 45;
      opCodes[4574] <= 45;
      opCodes[4658] <= 45;
      opCodes[4699] <= 45;
      opCodes[4740] <= 45;
      opCodes[4781] <= 45;
      opCodes[4822] <= 45;
      opCodes[4863] <= 45;
      opCodes[4904] <= 45;
      opCodes[4945] <= 45;
      opCodes[4965] <= 45;
      opCodes[4974] <= 45;
      opCodes[4993] <= 45;
      opCodes[5057] <= 45;
      opCodes[5098] <= 45;
      opCodes[5139] <= 45;
      opCodes[5180] <= 45;
      opCodes[5221] <= 45;
      opCodes[5262] <= 45;
      opCodes[5303] <= 45;
      opCodes[5344] <= 45;
      opCodes[5385] <= 45;
      opCodes[5490] <= 45;
      opCodes[5506] <= 45;
      opCodes[5546] <= 45;
      opCodes[5618] <= 45;
      opCodes[5656] <= 45;
      opCodes[5694] <= 45;
      opCodes[5732] <= 45;
      opCodes[5770] <= 45;
      opCodes[5802] <= 45;
      opCodes[5811] <= 45;
      opCodes[5814] <= 45;
      opCodes[5833] <= 45;
      opCodes[59] <= 46;
      opCodes[72] <= 46;
      opCodes[61] <= 47;
      opCodes[67] <= 48;
      opCodes[73] <= 49;
      opCodes[79] <= 50;
      opCodes[1253] <= 50;
      opCodes[1442] <= 50;
      opCodes[1781] <= 50;
      opCodes[80] <= 51;
      opCodes[86] <= 51;
      opCodes[110] <= 51;
      opCodes[123] <= 51;
      opCodes[1254] <= 51;
      opCodes[1260] <= 51;
      opCodes[1284] <= 51;
      opCodes[1297] <= 51;
      opCodes[1443] <= 51;
      opCodes[1449] <= 51;
      opCodes[1782] <= 51;
      opCodes[1788] <= 51;
      opCodes[1812] <= 51;
      opCodes[1825] <= 51;
      opCodes[5539] <= 51;
      opCodes[5554] <= 51;
      opCodes[5859] <= 51;
      opCodes[81] <= 52;
      opCodes[83] <= 52;
      opCodes[235] <= 52;
      opCodes[237] <= 52;
      opCodes[1255] <= 52;
      opCodes[1257] <= 52;
      opCodes[1444] <= 52;
      opCodes[1446] <= 52;
      opCodes[1783] <= 52;
      opCodes[1785] <= 52;
      opCodes[1972] <= 52;
      opCodes[1974] <= 52;
      opCodes[3603] <= 52;
      opCodes[3605] <= 52;
      opCodes[3665] <= 52;
      opCodes[3667] <= 52;
      opCodes[4602] <= 52;
      opCodes[4604] <= 52;
      opCodes[82] <= 53;
      opCodes[236] <= 53;
      opCodes[1256] <= 53;
      opCodes[1445] <= 53;
      opCodes[1784] <= 53;
      opCodes[1973] <= 53;
      opCodes[3604] <= 53;
      opCodes[3666] <= 53;
      opCodes[4603] <= 53;
      opCodes[84] <= 54;
      opCodes[238] <= 54;
      opCodes[1258] <= 54;
      opCodes[1447] <= 54;
      opCodes[1786] <= 54;
      opCodes[1975] <= 54;
      opCodes[3606] <= 54;
      opCodes[3668] <= 54;
      opCodes[4605] <= 54;
      opCodes[85] <= 55;
      opCodes[95] <= 56;
      opCodes[108] <= 56;
      opCodes[97] <= 57;
      opCodes[103] <= 58;
      opCodes[109] <= 59;
      opCodes[111] <= 60;
      opCodes[1285] <= 60;
      opCodes[1813] <= 60;
      opCodes[112] <= 61;
      opCodes[1286] <= 61;
      opCodes[1814] <= 61;
      opCodes[125] <= 62;
      opCodes[128] <= 62;
      opCodes[1299] <= 62;
      opCodes[1302] <= 62;
      opCodes[1827] <= 62;
      opCodes[1830] <= 62;
      opCodes[127] <= 63;
      opCodes[1301] <= 63;
      opCodes[1829] <= 63;
      opCodes[129] <= 64;
      opCodes[257] <= 64;
      opCodes[1303] <= 64;
      opCodes[1831] <= 64;
      opCodes[2744] <= 64;
      opCodes[4049] <= 64;
      opCodes[4986] <= 64;
      opCodes[5534] <= 64;
      opCodes[5549] <= 64;
      opCodes[5865] <= 64;
      opCodes[130] <= 65;
      opCodes[131] <= 66;
      opCodes[132] <= 67;
      opCodes[272] <= 67;
      opCodes[305] <= 67;
      opCodes[701] <= 67;
      opCodes[734] <= 67;
      opCodes[1306] <= 67;
      opCodes[1459] <= 67;
      opCodes[1834] <= 67;
      opCodes[5537] <= 67;
      opCodes[5564] <= 67;
      opCodes[5868] <= 67;
      opCodes[133] <= 68;
      opCodes[1307] <= 68;
      opCodes[1835] <= 68;
      opCodes[134] <= 69;
      opCodes[135] <= 70;
      opCodes[155] <= 70;
      opCodes[167] <= 70;
      opCodes[191] <= 70;
      opCodes[1309] <= 70;
      opCodes[1329] <= 70;
      opCodes[1341] <= 70;
      opCodes[1365] <= 70;
      opCodes[1837] <= 70;
      opCodes[1857] <= 70;
      opCodes[1869] <= 70;
      opCodes[1893] <= 70;
      opCodes[139] <= 71;
      opCodes[195] <= 71;
      opCodes[1313] <= 71;
      opCodes[1369] <= 71;
      opCodes[1841] <= 71;
      opCodes[1897] <= 71;
      opCodes[141] <= 72;
      opCodes[1315] <= 72;
      opCodes[1843] <= 72;
      opCodes[144] <= 73;
      opCodes[220] <= 73;
      opCodes[366] <= 73;
      opCodes[404] <= 73;
      opCodes[442] <= 73;
      opCodes[480] <= 73;
      opCodes[518] <= 73;
      opCodes[556] <= 73;
      opCodes[594] <= 73;
      opCodes[632] <= 73;
      opCodes[676] <= 73;
      opCodes[689] <= 73;
      opCodes[795] <= 73;
      opCodes[833] <= 73;
      opCodes[871] <= 73;
      opCodes[909] <= 73;
      opCodes[951] <= 73;
      opCodes[989] <= 73;
      opCodes[1027] <= 73;
      opCodes[1065] <= 73;
      opCodes[1103] <= 73;
      opCodes[1143] <= 73;
      opCodes[1159] <= 73;
      opCodes[1172] <= 73;
      opCodes[1318] <= 73;
      opCodes[1394] <= 73;
      opCodes[1520] <= 73;
      opCodes[1558] <= 73;
      opCodes[1596] <= 73;
      opCodes[1634] <= 73;
      opCodes[1700] <= 73;
      opCodes[1846] <= 73;
      opCodes[1922] <= 73;
      opCodes[2036] <= 73;
      opCodes[2077] <= 73;
      opCodes[2118] <= 73;
      opCodes[2159] <= 73;
      opCodes[2200] <= 73;
      opCodes[2241] <= 73;
      opCodes[2282] <= 73;
      opCodes[2323] <= 73;
      opCodes[2364] <= 73;
      opCodes[2405] <= 73;
      opCodes[2446] <= 73;
      opCodes[2487] <= 73;
      opCodes[2528] <= 73;
      opCodes[2569] <= 73;
      opCodes[2610] <= 73;
      opCodes[2651] <= 73;
      opCodes[2791] <= 73;
      opCodes[2832] <= 73;
      opCodes[2873] <= 73;
      opCodes[2914] <= 73;
      opCodes[2955] <= 73;
      opCodes[2996] <= 73;
      opCodes[3037] <= 73;
      opCodes[3078] <= 73;
      opCodes[3119] <= 73;
      opCodes[3143] <= 73;
      opCodes[3184] <= 73;
      opCodes[3225] <= 73;
      opCodes[3266] <= 73;
      opCodes[3307] <= 73;
      opCodes[3348] <= 73;
      opCodes[3389] <= 73;
      opCodes[3430] <= 73;
      opCodes[3471] <= 73;
      opCodes[3512] <= 73;
      opCodes[3536] <= 73;
      opCodes[3728] <= 73;
      opCodes[3769] <= 73;
      opCodes[3810] <= 73;
      opCodes[3851] <= 73;
      opCodes[3892] <= 73;
      opCodes[3933] <= 73;
      opCodes[3974] <= 73;
      opCodes[4015] <= 73;
      opCodes[4098] <= 73;
      opCodes[4162] <= 73;
      opCodes[4203] <= 73;
      opCodes[4244] <= 73;
      opCodes[4285] <= 73;
      opCodes[4326] <= 73;
      opCodes[4367] <= 73;
      opCodes[4408] <= 73;
      opCodes[4449] <= 73;
      opCodes[4490] <= 73;
      opCodes[4665] <= 73;
      opCodes[4706] <= 73;
      opCodes[4747] <= 73;
      opCodes[4788] <= 73;
      opCodes[4829] <= 73;
      opCodes[4870] <= 73;
      opCodes[4911] <= 73;
      opCodes[4952] <= 73;
      opCodes[5016] <= 73;
      opCodes[5064] <= 73;
      opCodes[5105] <= 73;
      opCodes[5146] <= 73;
      opCodes[5187] <= 73;
      opCodes[5228] <= 73;
      opCodes[5269] <= 73;
      opCodes[5310] <= 73;
      opCodes[5351] <= 73;
      opCodes[5392] <= 73;
      opCodes[5450] <= 73;
      opCodes[5625] <= 73;
      opCodes[5663] <= 73;
      opCodes[5701] <= 73;
      opCodes[5739] <= 73;
      opCodes[5781] <= 73;
      opCodes[5818] <= 73;
      opCodes[146] <= 74;
      opCodes[222] <= 74;
      opCodes[368] <= 74;
      opCodes[406] <= 74;
      opCodes[444] <= 74;
      opCodes[482] <= 74;
      opCodes[520] <= 74;
      opCodes[558] <= 74;
      opCodes[596] <= 74;
      opCodes[634] <= 74;
      opCodes[678] <= 74;
      opCodes[691] <= 74;
      opCodes[797] <= 74;
      opCodes[835] <= 74;
      opCodes[873] <= 74;
      opCodes[911] <= 74;
      opCodes[953] <= 74;
      opCodes[991] <= 74;
      opCodes[1029] <= 74;
      opCodes[1067] <= 74;
      opCodes[1105] <= 74;
      opCodes[1145] <= 74;
      opCodes[1161] <= 74;
      opCodes[1174] <= 74;
      opCodes[1320] <= 74;
      opCodes[1396] <= 74;
      opCodes[1522] <= 74;
      opCodes[1560] <= 74;
      opCodes[1598] <= 74;
      opCodes[1636] <= 74;
      opCodes[1702] <= 74;
      opCodes[1848] <= 74;
      opCodes[1924] <= 74;
      opCodes[2038] <= 74;
      opCodes[2079] <= 74;
      opCodes[2120] <= 74;
      opCodes[2161] <= 74;
      opCodes[2202] <= 74;
      opCodes[2243] <= 74;
      opCodes[2284] <= 74;
      opCodes[2325] <= 74;
      opCodes[2366] <= 74;
      opCodes[2407] <= 74;
      opCodes[2448] <= 74;
      opCodes[2489] <= 74;
      opCodes[2530] <= 74;
      opCodes[2571] <= 74;
      opCodes[2612] <= 74;
      opCodes[2653] <= 74;
      opCodes[2793] <= 74;
      opCodes[2834] <= 74;
      opCodes[2875] <= 74;
      opCodes[2916] <= 74;
      opCodes[2957] <= 74;
      opCodes[2998] <= 74;
      opCodes[3039] <= 74;
      opCodes[3080] <= 74;
      opCodes[3121] <= 74;
      opCodes[3145] <= 74;
      opCodes[3186] <= 74;
      opCodes[3227] <= 74;
      opCodes[3268] <= 74;
      opCodes[3309] <= 74;
      opCodes[3350] <= 74;
      opCodes[3391] <= 74;
      opCodes[3432] <= 74;
      opCodes[3473] <= 74;
      opCodes[3514] <= 74;
      opCodes[3538] <= 74;
      opCodes[3730] <= 74;
      opCodes[3771] <= 74;
      opCodes[3812] <= 74;
      opCodes[3853] <= 74;
      opCodes[3894] <= 74;
      opCodes[3935] <= 74;
      opCodes[3976] <= 74;
      opCodes[4017] <= 74;
      opCodes[4100] <= 74;
      opCodes[4164] <= 74;
      opCodes[4205] <= 74;
      opCodes[4246] <= 74;
      opCodes[4287] <= 74;
      opCodes[4328] <= 74;
      opCodes[4369] <= 74;
      opCodes[4410] <= 74;
      opCodes[4451] <= 74;
      opCodes[4492] <= 74;
      opCodes[4667] <= 74;
      opCodes[4708] <= 74;
      opCodes[4749] <= 74;
      opCodes[4790] <= 74;
      opCodes[4831] <= 74;
      opCodes[4872] <= 74;
      opCodes[4913] <= 74;
      opCodes[4954] <= 74;
      opCodes[5018] <= 74;
      opCodes[5066] <= 74;
      opCodes[5107] <= 74;
      opCodes[5148] <= 74;
      opCodes[5189] <= 74;
      opCodes[5230] <= 74;
      opCodes[5271] <= 74;
      opCodes[5312] <= 74;
      opCodes[5353] <= 74;
      opCodes[5394] <= 74;
      opCodes[5452] <= 74;
      opCodes[5627] <= 74;
      opCodes[5665] <= 74;
      opCodes[5703] <= 74;
      opCodes[5741] <= 74;
      opCodes[5783] <= 74;
      opCodes[5820] <= 74;
      opCodes[147] <= 75;
      opCodes[1321] <= 75;
      opCodes[1849] <= 75;
      opCodes[5019] <= 75;
      opCodes[5453] <= 75;
      opCodes[148] <= 76;
      opCodes[151] <= 77;
      opCodes[225] <= 77;
      opCodes[360] <= 77;
      opCodes[371] <= 77;
      opCodes[398] <= 77;
      opCodes[409] <= 77;
      opCodes[436] <= 77;
      opCodes[447] <= 77;
      opCodes[474] <= 77;
      opCodes[485] <= 77;
      opCodes[512] <= 77;
      opCodes[523] <= 77;
      opCodes[550] <= 77;
      opCodes[561] <= 77;
      opCodes[588] <= 77;
      opCodes[599] <= 77;
      opCodes[626] <= 77;
      opCodes[637] <= 77;
      opCodes[681] <= 77;
      opCodes[694] <= 77;
      opCodes[789] <= 77;
      opCodes[800] <= 77;
      opCodes[827] <= 77;
      opCodes[838] <= 77;
      opCodes[865] <= 77;
      opCodes[876] <= 77;
      opCodes[903] <= 77;
      opCodes[914] <= 77;
      opCodes[941] <= 77;
      opCodes[956] <= 77;
      opCodes[983] <= 77;
      opCodes[994] <= 77;
      opCodes[1021] <= 77;
      opCodes[1032] <= 77;
      opCodes[1059] <= 77;
      opCodes[1070] <= 77;
      opCodes[1097] <= 77;
      opCodes[1108] <= 77;
      opCodes[1135] <= 77;
      opCodes[1148] <= 77;
      opCodes[1164] <= 77;
      opCodes[1177] <= 77;
      opCodes[1325] <= 77;
      opCodes[1399] <= 77;
      opCodes[1514] <= 77;
      opCodes[1525] <= 77;
      opCodes[1552] <= 77;
      opCodes[1563] <= 77;
      opCodes[1590] <= 77;
      opCodes[1601] <= 77;
      opCodes[1628] <= 77;
      opCodes[1639] <= 77;
      opCodes[1705] <= 77;
      opCodes[1853] <= 77;
      opCodes[1927] <= 77;
      opCodes[2030] <= 77;
      opCodes[2041] <= 77;
      opCodes[2071] <= 77;
      opCodes[2082] <= 77;
      opCodes[2112] <= 77;
      opCodes[2123] <= 77;
      opCodes[2153] <= 77;
      opCodes[2164] <= 77;
      opCodes[2194] <= 77;
      opCodes[2205] <= 77;
      opCodes[2235] <= 77;
      opCodes[2246] <= 77;
      opCodes[2276] <= 77;
      opCodes[2287] <= 77;
      opCodes[2317] <= 77;
      opCodes[2328] <= 77;
      opCodes[2358] <= 77;
      opCodes[2369] <= 77;
      opCodes[2399] <= 77;
      opCodes[2410] <= 77;
      opCodes[2440] <= 77;
      opCodes[2451] <= 77;
      opCodes[2481] <= 77;
      opCodes[2492] <= 77;
      opCodes[2522] <= 77;
      opCodes[2533] <= 77;
      opCodes[2563] <= 77;
      opCodes[2574] <= 77;
      opCodes[2604] <= 77;
      opCodes[2615] <= 77;
      opCodes[2645] <= 77;
      opCodes[2656] <= 77;
      opCodes[2785] <= 77;
      opCodes[2796] <= 77;
      opCodes[2826] <= 77;
      opCodes[2837] <= 77;
      opCodes[2867] <= 77;
      opCodes[2878] <= 77;
      opCodes[2908] <= 77;
      opCodes[2919] <= 77;
      opCodes[2949] <= 77;
      opCodes[2960] <= 77;
      opCodes[2990] <= 77;
      opCodes[3001] <= 77;
      opCodes[3031] <= 77;
      opCodes[3042] <= 77;
      opCodes[3072] <= 77;
      opCodes[3083] <= 77;
      opCodes[3113] <= 77;
      opCodes[3124] <= 77;
      opCodes[3148] <= 77;
      opCodes[3178] <= 77;
      opCodes[3189] <= 77;
      opCodes[3219] <= 77;
      opCodes[3230] <= 77;
      opCodes[3260] <= 77;
      opCodes[3271] <= 77;
      opCodes[3301] <= 77;
      opCodes[3312] <= 77;
      opCodes[3342] <= 77;
      opCodes[3353] <= 77;
      opCodes[3383] <= 77;
      opCodes[3394] <= 77;
      opCodes[3424] <= 77;
      opCodes[3435] <= 77;
      opCodes[3465] <= 77;
      opCodes[3476] <= 77;
      opCodes[3506] <= 77;
      opCodes[3517] <= 77;
      opCodes[3541] <= 77;
      opCodes[3700] <= 77;
      opCodes[3733] <= 77;
      opCodes[3741] <= 77;
      opCodes[3774] <= 77;
      opCodes[3782] <= 77;
      opCodes[3815] <= 77;
      opCodes[3823] <= 77;
      opCodes[3856] <= 77;
      opCodes[3864] <= 77;
      opCodes[3897] <= 77;
      opCodes[3905] <= 77;
      opCodes[3938] <= 77;
      opCodes[3946] <= 77;
      opCodes[3979] <= 77;
      opCodes[3987] <= 77;
      opCodes[4020] <= 77;
      opCodes[4103] <= 77;
      opCodes[4108] <= 77;
      opCodes[4134] <= 77;
      opCodes[4167] <= 77;
      opCodes[4175] <= 77;
      opCodes[4208] <= 77;
      opCodes[4216] <= 77;
      opCodes[4249] <= 77;
      opCodes[4257] <= 77;
      opCodes[4290] <= 77;
      opCodes[4298] <= 77;
      opCodes[4331] <= 77;
      opCodes[4339] <= 77;
      opCodes[4372] <= 77;
      opCodes[4380] <= 77;
      opCodes[4413] <= 77;
      opCodes[4421] <= 77;
      opCodes[4454] <= 77;
      opCodes[4462] <= 77;
      opCodes[4495] <= 77;
      opCodes[4559] <= 77;
      opCodes[4659] <= 77;
      opCodes[4670] <= 77;
      opCodes[4700] <= 77;
      opCodes[4711] <= 77;
      opCodes[4741] <= 77;
      opCodes[4752] <= 77;
      opCodes[4782] <= 77;
      opCodes[4793] <= 77;
      opCodes[4823] <= 77;
      opCodes[4834] <= 77;
      opCodes[4864] <= 77;
      opCodes[4875] <= 77;
      opCodes[4905] <= 77;
      opCodes[4916] <= 77;
      opCodes[4946] <= 77;
      opCodes[4957] <= 77;
      opCodes[5023] <= 77;
      opCodes[5058] <= 77;
      opCodes[5069] <= 77;
      opCodes[5099] <= 77;
      opCodes[5110] <= 77;
      opCodes[5140] <= 77;
      opCodes[5151] <= 77;
      opCodes[5181] <= 77;
      opCodes[5192] <= 77;
      opCodes[5222] <= 77;
      opCodes[5233] <= 77;
      opCodes[5263] <= 77;
      opCodes[5274] <= 77;
      opCodes[5304] <= 77;
      opCodes[5315] <= 77;
      opCodes[5345] <= 77;
      opCodes[5356] <= 77;
      opCodes[5386] <= 77;
      opCodes[5397] <= 77;
      opCodes[5457] <= 77;
      opCodes[5491] <= 77;
      opCodes[5619] <= 77;
      opCodes[5630] <= 77;
      opCodes[5657] <= 77;
      opCodes[5668] <= 77;
      opCodes[5695] <= 77;
      opCodes[5706] <= 77;
      opCodes[5733] <= 77;
      opCodes[5744] <= 77;
      opCodes[5771] <= 77;
      opCodes[5786] <= 77;
      opCodes[5823] <= 77;
      opCodes[152] <= 78;
      opCodes[226] <= 78;
      opCodes[1326] <= 78;
      opCodes[1400] <= 78;
      opCodes[1854] <= 78;
      opCodes[1928] <= 78;
      opCodes[153] <= 79;
      opCodes[227] <= 79;
      opCodes[230] <= 79;
      opCodes[1327] <= 79;
      opCodes[1401] <= 79;
      opCodes[1404] <= 79;
      opCodes[1855] <= 79;
      opCodes[1929] <= 79;
      opCodes[1932] <= 79;
      opCodes[154] <= 80;
      opCodes[228] <= 80;
      opCodes[156] <= 81;
      opCodes[164] <= 81;
      opCodes[247] <= 81;
      opCodes[259] <= 81;
      opCodes[1330] <= 81;
      opCodes[1338] <= 81;
      opCodes[1858] <= 81;
      opCodes[1866] <= 81;
      opCodes[5540] <= 81;
      opCodes[5551] <= 81;
      opCodes[157] <= 82;
      opCodes[165] <= 82;
      opCodes[234] <= 82;
      opCodes[240] <= 82;
      opCodes[249] <= 82;
      opCodes[260] <= 82;
      opCodes[1331] <= 82;
      opCodes[1339] <= 82;
      opCodes[1859] <= 82;
      opCodes[1867] <= 82;
      opCodes[5541] <= 82;
      opCodes[5552] <= 82;
      opCodes[5857] <= 82;
      opCodes[158] <= 83;
      opCodes[160] <= 83;
      opCodes[241] <= 83;
      opCodes[243] <= 83;
      opCodes[1332] <= 83;
      opCodes[1334] <= 83;
      opCodes[1860] <= 83;
      opCodes[1862] <= 83;
      opCodes[1980] <= 83;
      opCodes[1982] <= 83;
      opCodes[1986] <= 83;
      opCodes[1988] <= 83;
      opCodes[3673] <= 83;
      opCodes[3675] <= 83;
      opCodes[3679] <= 83;
      opCodes[3681] <= 83;
      opCodes[4610] <= 83;
      opCodes[4612] <= 83;
      opCodes[4616] <= 83;
      opCodes[4618] <= 83;
      opCodes[159] <= 84;
      opCodes[242] <= 84;
      opCodes[1333] <= 84;
      opCodes[1861] <= 84;
      opCodes[1981] <= 84;
      opCodes[1987] <= 84;
      opCodes[3674] <= 84;
      opCodes[3680] <= 84;
      opCodes[4611] <= 84;
      opCodes[4617] <= 84;
      opCodes[161] <= 85;
      opCodes[244] <= 85;
      opCodes[1335] <= 85;
      opCodes[1863] <= 85;
      opCodes[1983] <= 85;
      opCodes[1989] <= 85;
      opCodes[3676] <= 85;
      opCodes[3682] <= 85;
      opCodes[4613] <= 85;
      opCodes[4619] <= 85;
      opCodes[162] <= 86;
      opCodes[245] <= 86;
      opCodes[1336] <= 86;
      opCodes[1864] <= 86;
      opCodes[1996] <= 86;
      opCodes[3085] <= 86;
      opCodes[3478] <= 86;
      opCodes[3689] <= 86;
      opCodes[4456] <= 86;
      opCodes[4626] <= 86;
      opCodes[5358] <= 86;
      opCodes[163] <= 87;
      opCodes[246] <= 87;
      opCodes[258] <= 87;
      opCodes[1337] <= 87;
      opCodes[1865] <= 87;
      opCodes[5550] <= 87;
      opCodes[166] <= 88;
      opCodes[176] <= 89;
      opCodes[189] <= 89;
      opCodes[178] <= 90;
      opCodes[184] <= 91;
      opCodes[190] <= 92;
      opCodes[198] <= 93;
      opCodes[1372] <= 93;
      opCodes[1678] <= 93;
      opCodes[1900] <= 93;
      opCodes[5796] <= 93;
      opCodes[200] <= 94;
      opCodes[214] <= 94;
      opCodes[1374] <= 94;
      opCodes[1388] <= 94;
      opCodes[1680] <= 94;
      opCodes[1694] <= 94;
      opCodes[1902] <= 94;
      opCodes[1916] <= 94;
      opCodes[5798] <= 94;
      opCodes[5812] <= 94;
      opCodes[201] <= 95;
      opCodes[212] <= 95;
      opCodes[1375] <= 95;
      opCodes[1386] <= 95;
      opCodes[1681] <= 95;
      opCodes[1692] <= 95;
      opCodes[1903] <= 95;
      opCodes[1914] <= 95;
      opCodes[5799] <= 95;
      opCodes[5810] <= 95;
      opCodes[202] <= 96;
      opCodes[205] <= 96;
      opCodes[217] <= 96;
      opCodes[1376] <= 96;
      opCodes[1379] <= 96;
      opCodes[1391] <= 96;
      opCodes[1682] <= 96;
      opCodes[1685] <= 96;
      opCodes[1697] <= 96;
      opCodes[1904] <= 96;
      opCodes[1907] <= 96;
      opCodes[1919] <= 96;
      opCodes[5800] <= 96;
      opCodes[5803] <= 96;
      opCodes[5815] <= 96;
      opCodes[203] <= 97;
      opCodes[215] <= 97;
      opCodes[1377] <= 97;
      opCodes[1389] <= 97;
      opCodes[1683] <= 97;
      opCodes[1695] <= 97;
      opCodes[1905] <= 97;
      opCodes[1917] <= 97;
      opCodes[5801] <= 97;
      opCodes[5813] <= 97;
      opCodes[206] <= 98;
      opCodes[1380] <= 98;
      opCodes[1686] <= 98;
      opCodes[1908] <= 98;
      opCodes[5804] <= 98;
      opCodes[207] <= 99;
      opCodes[208] <= 100;
      opCodes[1382] <= 100;
      opCodes[1688] <= 100;
      opCodes[1910] <= 100;
      opCodes[5806] <= 100;
      opCodes[209] <= 101;
      opCodes[1383] <= 101;
      opCodes[1689] <= 101;
      opCodes[1911] <= 101;
      opCodes[5807] <= 101;
      opCodes[210] <= 102;
      opCodes[1384] <= 102;
      opCodes[1690] <= 102;
      opCodes[1912] <= 102;
      opCodes[5808] <= 102;
      opCodes[211] <= 103;
      opCodes[1385] <= 103;
      opCodes[1691] <= 103;
      opCodes[1913] <= 103;
      opCodes[5809] <= 103;
      opCodes[218] <= 104;
      opCodes[229] <= 105;
      opCodes[1403] <= 105;
      opCodes[1931] <= 105;
      opCodes[231] <= 106;
      opCodes[1405] <= 106;
      opCodes[232] <= 107;
      opCodes[1406] <= 107;
      opCodes[233] <= 108;
      opCodes[239] <= 109;
      opCodes[248] <= 110;
      opCodes[250] <= 111;
      opCodes[252] <= 111;
      opCodes[255] <= 111;
      opCodes[1941] <= 111;
      opCodes[1944] <= 111;
      opCodes[2719] <= 111;
      opCodes[2721] <= 111;
      opCodes[2724] <= 111;
      opCodes[2728] <= 111;
      opCodes[2730] <= 111;
      opCodes[2733] <= 111;
      opCodes[3609] <= 111;
      opCodes[3611] <= 111;
      opCodes[3614] <= 111;
      opCodes[3631] <= 111;
      opCodes[3633] <= 111;
      opCodes[3636] <= 111;
      opCodes[4024] <= 111;
      opCodes[4026] <= 111;
      opCodes[4029] <= 111;
      opCodes[4033] <= 111;
      opCodes[4035] <= 111;
      opCodes[4038] <= 111;
      opCodes[4116] <= 111;
      opCodes[4118] <= 111;
      opCodes[4121] <= 111;
      opCodes[4961] <= 111;
      opCodes[4963] <= 111;
      opCodes[4966] <= 111;
      opCodes[4970] <= 111;
      opCodes[4972] <= 111;
      opCodes[4975] <= 111;
      opCodes[5542] <= 111;
      opCodes[5544] <= 111;
      opCodes[5547] <= 111;
      opCodes[251] <= 112;
      opCodes[1940] <= 112;
      opCodes[2720] <= 112;
      opCodes[2729] <= 112;
      opCodes[3610] <= 112;
      opCodes[3632] <= 112;
      opCodes[4025] <= 112;
      opCodes[4034] <= 112;
      opCodes[4117] <= 112;
      opCodes[4962] <= 112;
      opCodes[4971] <= 112;
      opCodes[5543] <= 112;
      opCodes[253] <= 113;
      opCodes[256] <= 113;
      opCodes[1942] <= 113;
      opCodes[1945] <= 113;
      opCodes[2722] <= 113;
      opCodes[2725] <= 113;
      opCodes[2731] <= 113;
      opCodes[2734] <= 113;
      opCodes[3612] <= 113;
      opCodes[3615] <= 113;
      opCodes[3634] <= 113;
      opCodes[3637] <= 113;
      opCodes[4027] <= 113;
      opCodes[4030] <= 113;
      opCodes[4036] <= 113;
      opCodes[4039] <= 113;
      opCodes[4119] <= 113;
      opCodes[4122] <= 113;
      opCodes[4964] <= 113;
      opCodes[4967] <= 113;
      opCodes[4973] <= 113;
      opCodes[4976] <= 113;
      opCodes[5545] <= 113;
      opCodes[5548] <= 113;
      opCodes[261] <= 114;
      opCodes[262] <= 115;
      opCodes[263] <= 116;
      opCodes[267] <= 117;
      opCodes[268] <= 118;
      opCodes[301] <= 118;
      opCodes[697] <= 118;
      opCodes[730] <= 118;
      opCodes[1455] <= 118;
      opCodes[2684] <= 118;
      opCodes[2712] <= 118;
      opCodes[3566] <= 118;
      opCodes[3594] <= 118;
      opCodes[4520] <= 118;
      opCodes[5422] <= 118;
      opCodes[5560] <= 118;
      opCodes[269] <= 119;
      opCodes[270] <= 120;
      opCodes[298] <= 120;
      opCodes[361] <= 120;
      opCodes[399] <= 120;
      opCodes[437] <= 120;
      opCodes[475] <= 120;
      opCodes[645] <= 120;
      opCodes[671] <= 120;
      opCodes[271] <= 121;
      opCodes[273] <= 122;
      opCodes[274] <= 123;
      opCodes[307] <= 123;
      opCodes[703] <= 123;
      opCodes[736] <= 123;
      opCodes[1461] <= 123;
      opCodes[2687] <= 123;
      opCodes[2715] <= 123;
      opCodes[3569] <= 123;
      opCodes[3597] <= 123;
      opCodes[4523] <= 123;
      opCodes[5425] <= 123;
      opCodes[5566] <= 123;
      opCodes[275] <= 124;
      opCodes[276] <= 125;
      opCodes[277] <= 126;
      opCodes[278] <= 127;
      opCodes[311] <= 127;
      opCodes[707] <= 127;
      opCodes[740] <= 127;
      opCodes[1465] <= 127;
      opCodes[5570] <= 127;
      opCodes[279] <= 128;
      opCodes[312] <= 128;
      opCodes[708] <= 128;
      opCodes[741] <= 128;
      opCodes[1466] <= 128;
      opCodes[5571] <= 128;
      opCodes[280] <= 129;
      opCodes[313] <= 129;
      opCodes[709] <= 129;
      opCodes[742] <= 129;
      opCodes[1467] <= 129;
      opCodes[5572] <= 129;
      opCodes[281] <= 130;
      opCodes[314] <= 130;
      opCodes[710] <= 130;
      opCodes[743] <= 130;
      opCodes[1468] <= 130;
      opCodes[5573] <= 130;
      opCodes[282] <= 131;
      opCodes[315] <= 131;
      opCodes[711] <= 131;
      opCodes[744] <= 131;
      opCodes[1469] <= 131;
      opCodes[5574] <= 131;
      opCodes[283] <= 132;
      opCodes[316] <= 132;
      opCodes[712] <= 132;
      opCodes[745] <= 132;
      opCodes[1470] <= 132;
      opCodes[5575] <= 132;
      opCodes[284] <= 133;
      opCodes[317] <= 133;
      opCodes[713] <= 133;
      opCodes[746] <= 133;
      opCodes[1471] <= 133;
      opCodes[5576] <= 133;
      opCodes[285] <= 134;
      opCodes[318] <= 134;
      opCodes[714] <= 134;
      opCodes[747] <= 134;
      opCodes[1472] <= 134;
      opCodes[5577] <= 134;
      opCodes[286] <= 135;
      opCodes[319] <= 135;
      opCodes[715] <= 135;
      opCodes[748] <= 135;
      opCodes[1473] <= 135;
      opCodes[5578] <= 135;
      opCodes[287] <= 136;
      opCodes[320] <= 136;
      opCodes[716] <= 136;
      opCodes[749] <= 136;
      opCodes[1474] <= 136;
      opCodes[5579] <= 136;
      opCodes[288] <= 137;
      opCodes[321] <= 137;
      opCodes[717] <= 137;
      opCodes[750] <= 137;
      opCodes[1475] <= 137;
      opCodes[5580] <= 137;
      opCodes[289] <= 138;
      opCodes[322] <= 138;
      opCodes[718] <= 138;
      opCodes[751] <= 138;
      opCodes[1476] <= 138;
      opCodes[5581] <= 138;
      opCodes[290] <= 139;
      opCodes[323] <= 139;
      opCodes[719] <= 139;
      opCodes[752] <= 139;
      opCodes[1477] <= 139;
      opCodes[5582] <= 139;
      opCodes[291] <= 140;
      opCodes[324] <= 140;
      opCodes[720] <= 140;
      opCodes[753] <= 140;
      opCodes[1478] <= 140;
      opCodes[5583] <= 140;
      opCodes[292] <= 141;
      opCodes[325] <= 141;
      opCodes[721] <= 141;
      opCodes[754] <= 141;
      opCodes[1479] <= 141;
      opCodes[5584] <= 141;
      opCodes[293] <= 142;
      opCodes[326] <= 142;
      opCodes[722] <= 142;
      opCodes[755] <= 142;
      opCodes[1480] <= 142;
      opCodes[5585] <= 142;
      opCodes[294] <= 143;
      opCodes[327] <= 143;
      opCodes[723] <= 143;
      opCodes[756] <= 143;
      opCodes[1481] <= 143;
      opCodes[5586] <= 143;
      opCodes[295] <= 144;
      opCodes[328] <= 144;
      opCodes[724] <= 144;
      opCodes[757] <= 144;
      opCodes[1482] <= 144;
      opCodes[5587] <= 144;
      opCodes[296] <= 145;
      opCodes[329] <= 145;
      opCodes[725] <= 145;
      opCodes[758] <= 145;
      opCodes[1483] <= 145;
      opCodes[5588] <= 145;
      opCodes[297] <= 146;
      opCodes[330] <= 146;
      opCodes[726] <= 146;
      opCodes[759] <= 146;
      opCodes[1484] <= 146;
      opCodes[5589] <= 146;
      opCodes[299] <= 147;
      opCodes[332] <= 147;
      opCodes[1486] <= 147;
      opCodes[2658] <= 147;
      opCodes[300] <= 148;
      opCodes[333] <= 148;
      opCodes[1487] <= 148;
      opCodes[2659] <= 148;
      opCodes[302] <= 149;
      opCodes[303] <= 150;
      opCodes[331] <= 150;
      opCodes[513] <= 150;
      opCodes[551] <= 150;
      opCodes[589] <= 150;
      opCodes[627] <= 150;
      opCodes[684] <= 150;
      opCodes[304] <= 151;
      opCodes[306] <= 152;
      opCodes[308] <= 153;
      opCodes[309] <= 154;
      opCodes[310] <= 155;
      opCodes[336] <= 156;
      opCodes[374] <= 156;
      opCodes[412] <= 156;
      opCodes[450] <= 156;
      opCodes[488] <= 156;
      opCodes[526] <= 156;
      opCodes[564] <= 156;
      opCodes[602] <= 156;
      opCodes[765] <= 156;
      opCodes[803] <= 156;
      opCodes[841] <= 156;
      opCodes[879] <= 156;
      opCodes[917] <= 156;
      opCodes[959] <= 156;
      opCodes[997] <= 156;
      opCodes[1035] <= 156;
      opCodes[1073] <= 156;
      opCodes[1111] <= 156;
      opCodes[1490] <= 156;
      opCodes[1528] <= 156;
      opCodes[1566] <= 156;
      opCodes[1604] <= 156;
      opCodes[2006] <= 156;
      opCodes[2047] <= 156;
      opCodes[2088] <= 156;
      opCodes[2129] <= 156;
      opCodes[2170] <= 156;
      opCodes[2211] <= 156;
      opCodes[2252] <= 156;
      opCodes[2293] <= 156;
      opCodes[2334] <= 156;
      opCodes[2375] <= 156;
      opCodes[2416] <= 156;
      opCodes[2457] <= 156;
      opCodes[2498] <= 156;
      opCodes[2539] <= 156;
      opCodes[2580] <= 156;
      opCodes[2621] <= 156;
      opCodes[2761] <= 156;
      opCodes[2802] <= 156;
      opCodes[2843] <= 156;
      opCodes[2884] <= 156;
      opCodes[2925] <= 156;
      opCodes[2966] <= 156;
      opCodes[3007] <= 156;
      opCodes[3048] <= 156;
      opCodes[3089] <= 156;
      opCodes[3154] <= 156;
      opCodes[3195] <= 156;
      opCodes[3236] <= 156;
      opCodes[3277] <= 156;
      opCodes[3318] <= 156;
      opCodes[3359] <= 156;
      opCodes[3400] <= 156;
      opCodes[3441] <= 156;
      opCodes[3482] <= 156;
      opCodes[4635] <= 156;
      opCodes[4676] <= 156;
      opCodes[4717] <= 156;
      opCodes[4758] <= 156;
      opCodes[4799] <= 156;
      opCodes[4840] <= 156;
      opCodes[4881] <= 156;
      opCodes[4922] <= 156;
      opCodes[5034] <= 156;
      opCodes[5075] <= 156;
      opCodes[5116] <= 156;
      opCodes[5157] <= 156;
      opCodes[5198] <= 156;
      opCodes[5239] <= 156;
      opCodes[5280] <= 156;
      opCodes[5321] <= 156;
      opCodes[5362] <= 156;
      opCodes[5595] <= 156;
      opCodes[5633] <= 156;
      opCodes[5671] <= 156;
      opCodes[5709] <= 156;
      opCodes[5747] <= 156;
      opCodes[342] <= 157;
      opCodes[380] <= 157;
      opCodes[418] <= 157;
      opCodes[456] <= 157;
      opCodes[494] <= 157;
      opCodes[532] <= 157;
      opCodes[570] <= 157;
      opCodes[608] <= 157;
      opCodes[771] <= 157;
      opCodes[809] <= 157;
      opCodes[847] <= 157;
      opCodes[885] <= 157;
      opCodes[923] <= 157;
      opCodes[965] <= 157;
      opCodes[1003] <= 157;
      opCodes[1041] <= 157;
      opCodes[1079] <= 157;
      opCodes[1117] <= 157;
      opCodes[1496] <= 157;
      opCodes[1534] <= 157;
      opCodes[1572] <= 157;
      opCodes[1610] <= 157;
      opCodes[2012] <= 157;
      opCodes[2053] <= 157;
      opCodes[2094] <= 157;
      opCodes[2135] <= 157;
      opCodes[2176] <= 157;
      opCodes[2217] <= 157;
      opCodes[2258] <= 157;
      opCodes[2299] <= 157;
      opCodes[2340] <= 157;
      opCodes[2381] <= 157;
      opCodes[2422] <= 157;
      opCodes[2463] <= 157;
      opCodes[2504] <= 157;
      opCodes[2545] <= 157;
      opCodes[2586] <= 157;
      opCodes[2627] <= 157;
      opCodes[2767] <= 157;
      opCodes[2808] <= 157;
      opCodes[2849] <= 157;
      opCodes[2890] <= 157;
      opCodes[2931] <= 157;
      opCodes[2972] <= 157;
      opCodes[3013] <= 157;
      opCodes[3054] <= 157;
      opCodes[3095] <= 157;
      opCodes[3160] <= 157;
      opCodes[3201] <= 157;
      opCodes[3242] <= 157;
      opCodes[3283] <= 157;
      opCodes[3324] <= 157;
      opCodes[3365] <= 157;
      opCodes[3406] <= 157;
      opCodes[3447] <= 157;
      opCodes[3488] <= 157;
      opCodes[4641] <= 157;
      opCodes[4682] <= 157;
      opCodes[4723] <= 157;
      opCodes[4764] <= 157;
      opCodes[4805] <= 157;
      opCodes[4846] <= 157;
      opCodes[4887] <= 157;
      opCodes[4928] <= 157;
      opCodes[5040] <= 157;
      opCodes[5081] <= 157;
      opCodes[5122] <= 157;
      opCodes[5163] <= 157;
      opCodes[5204] <= 157;
      opCodes[5245] <= 157;
      opCodes[5286] <= 157;
      opCodes[5327] <= 157;
      opCodes[5368] <= 157;
      opCodes[5601] <= 157;
      opCodes[5639] <= 157;
      opCodes[5677] <= 157;
      opCodes[5715] <= 157;
      opCodes[5753] <= 157;
      opCodes[343] <= 158;
      opCodes[381] <= 158;
      opCodes[419] <= 158;
      opCodes[457] <= 158;
      opCodes[495] <= 158;
      opCodes[533] <= 158;
      opCodes[571] <= 158;
      opCodes[609] <= 158;
      opCodes[772] <= 158;
      opCodes[810] <= 158;
      opCodes[848] <= 158;
      opCodes[886] <= 158;
      opCodes[924] <= 158;
      opCodes[966] <= 158;
      opCodes[1004] <= 158;
      opCodes[1042] <= 158;
      opCodes[1080] <= 158;
      opCodes[1118] <= 158;
      opCodes[1497] <= 158;
      opCodes[1535] <= 158;
      opCodes[1573] <= 158;
      opCodes[1611] <= 158;
      opCodes[2013] <= 158;
      opCodes[2054] <= 158;
      opCodes[2095] <= 158;
      opCodes[2136] <= 158;
      opCodes[2177] <= 158;
      opCodes[2218] <= 158;
      opCodes[2259] <= 158;
      opCodes[2300] <= 158;
      opCodes[2341] <= 158;
      opCodes[2382] <= 158;
      opCodes[2423] <= 158;
      opCodes[2464] <= 158;
      opCodes[2505] <= 158;
      opCodes[2546] <= 158;
      opCodes[2587] <= 158;
      opCodes[2628] <= 158;
      opCodes[2768] <= 158;
      opCodes[2809] <= 158;
      opCodes[2850] <= 158;
      opCodes[2891] <= 158;
      opCodes[2932] <= 158;
      opCodes[2973] <= 158;
      opCodes[3014] <= 158;
      opCodes[3055] <= 158;
      opCodes[3096] <= 158;
      opCodes[3161] <= 158;
      opCodes[3202] <= 158;
      opCodes[3243] <= 158;
      opCodes[3284] <= 158;
      opCodes[3325] <= 158;
      opCodes[3366] <= 158;
      opCodes[3407] <= 158;
      opCodes[3448] <= 158;
      opCodes[3489] <= 158;
      opCodes[4642] <= 158;
      opCodes[4683] <= 158;
      opCodes[4724] <= 158;
      opCodes[4765] <= 158;
      opCodes[4806] <= 158;
      opCodes[4847] <= 158;
      opCodes[4888] <= 158;
      opCodes[4929] <= 158;
      opCodes[5041] <= 158;
      opCodes[5082] <= 158;
      opCodes[5123] <= 158;
      opCodes[5164] <= 158;
      opCodes[5205] <= 158;
      opCodes[5246] <= 158;
      opCodes[5287] <= 158;
      opCodes[5328] <= 158;
      opCodes[5369] <= 158;
      opCodes[5602] <= 158;
      opCodes[5640] <= 158;
      opCodes[5678] <= 158;
      opCodes[5716] <= 158;
      opCodes[5754] <= 158;
      opCodes[344] <= 159;
      opCodes[382] <= 159;
      opCodes[420] <= 159;
      opCodes[458] <= 159;
      opCodes[496] <= 159;
      opCodes[534] <= 159;
      opCodes[572] <= 159;
      opCodes[610] <= 159;
      opCodes[773] <= 159;
      opCodes[811] <= 159;
      opCodes[849] <= 159;
      opCodes[887] <= 159;
      opCodes[925] <= 159;
      opCodes[967] <= 159;
      opCodes[1005] <= 159;
      opCodes[1043] <= 159;
      opCodes[1081] <= 159;
      opCodes[1119] <= 159;
      opCodes[1498] <= 159;
      opCodes[1536] <= 159;
      opCodes[1574] <= 159;
      opCodes[1612] <= 159;
      opCodes[2014] <= 159;
      opCodes[2055] <= 159;
      opCodes[2096] <= 159;
      opCodes[2137] <= 159;
      opCodes[2178] <= 159;
      opCodes[2219] <= 159;
      opCodes[2260] <= 159;
      opCodes[2301] <= 159;
      opCodes[2342] <= 159;
      opCodes[2383] <= 159;
      opCodes[2424] <= 159;
      opCodes[2465] <= 159;
      opCodes[2506] <= 159;
      opCodes[2547] <= 159;
      opCodes[2588] <= 159;
      opCodes[2629] <= 159;
      opCodes[2769] <= 159;
      opCodes[2810] <= 159;
      opCodes[2851] <= 159;
      opCodes[2892] <= 159;
      opCodes[2933] <= 159;
      opCodes[2974] <= 159;
      opCodes[3015] <= 159;
      opCodes[3056] <= 159;
      opCodes[3097] <= 159;
      opCodes[3162] <= 159;
      opCodes[3203] <= 159;
      opCodes[3244] <= 159;
      opCodes[3285] <= 159;
      opCodes[3326] <= 159;
      opCodes[3367] <= 159;
      opCodes[3408] <= 159;
      opCodes[3449] <= 159;
      opCodes[3490] <= 159;
      opCodes[4643] <= 159;
      opCodes[4684] <= 159;
      opCodes[4725] <= 159;
      opCodes[4766] <= 159;
      opCodes[4807] <= 159;
      opCodes[4848] <= 159;
      opCodes[4889] <= 159;
      opCodes[4930] <= 159;
      opCodes[5042] <= 159;
      opCodes[5083] <= 159;
      opCodes[5124] <= 159;
      opCodes[5165] <= 159;
      opCodes[5206] <= 159;
      opCodes[5247] <= 159;
      opCodes[5288] <= 159;
      opCodes[5329] <= 159;
      opCodes[5370] <= 159;
      opCodes[5603] <= 159;
      opCodes[5641] <= 159;
      opCodes[5679] <= 159;
      opCodes[5717] <= 159;
      opCodes[5755] <= 159;
      opCodes[345] <= 160;
      opCodes[383] <= 160;
      opCodes[421] <= 160;
      opCodes[459] <= 160;
      opCodes[497] <= 160;
      opCodes[535] <= 160;
      opCodes[573] <= 160;
      opCodes[611] <= 160;
      opCodes[774] <= 160;
      opCodes[812] <= 160;
      opCodes[850] <= 160;
      opCodes[888] <= 160;
      opCodes[926] <= 160;
      opCodes[968] <= 160;
      opCodes[1006] <= 160;
      opCodes[1044] <= 160;
      opCodes[1082] <= 160;
      opCodes[1120] <= 160;
      opCodes[1499] <= 160;
      opCodes[1537] <= 160;
      opCodes[1575] <= 160;
      opCodes[1613] <= 160;
      opCodes[2015] <= 160;
      opCodes[2056] <= 160;
      opCodes[2097] <= 160;
      opCodes[2138] <= 160;
      opCodes[2179] <= 160;
      opCodes[2220] <= 160;
      opCodes[2261] <= 160;
      opCodes[2302] <= 160;
      opCodes[2343] <= 160;
      opCodes[2384] <= 160;
      opCodes[2425] <= 160;
      opCodes[2466] <= 160;
      opCodes[2507] <= 160;
      opCodes[2548] <= 160;
      opCodes[2589] <= 160;
      opCodes[2630] <= 160;
      opCodes[2770] <= 160;
      opCodes[2811] <= 160;
      opCodes[2852] <= 160;
      opCodes[2893] <= 160;
      opCodes[2934] <= 160;
      opCodes[2975] <= 160;
      opCodes[3016] <= 160;
      opCodes[3057] <= 160;
      opCodes[3098] <= 160;
      opCodes[3163] <= 160;
      opCodes[3204] <= 160;
      opCodes[3245] <= 160;
      opCodes[3286] <= 160;
      opCodes[3327] <= 160;
      opCodes[3368] <= 160;
      opCodes[3409] <= 160;
      opCodes[3450] <= 160;
      opCodes[3491] <= 160;
      opCodes[4644] <= 160;
      opCodes[4685] <= 160;
      opCodes[4726] <= 160;
      opCodes[4767] <= 160;
      opCodes[4808] <= 160;
      opCodes[4849] <= 160;
      opCodes[4890] <= 160;
      opCodes[4931] <= 160;
      opCodes[5043] <= 160;
      opCodes[5084] <= 160;
      opCodes[5125] <= 160;
      opCodes[5166] <= 160;
      opCodes[5207] <= 160;
      opCodes[5248] <= 160;
      opCodes[5289] <= 160;
      opCodes[5330] <= 160;
      opCodes[5371] <= 160;
      opCodes[5604] <= 160;
      opCodes[5642] <= 160;
      opCodes[5680] <= 160;
      opCodes[5718] <= 160;
      opCodes[5756] <= 160;
      opCodes[346] <= 161;
      opCodes[347] <= 162;
      opCodes[385] <= 162;
      opCodes[423] <= 162;
      opCodes[461] <= 162;
      opCodes[499] <= 162;
      opCodes[537] <= 162;
      opCodes[575] <= 162;
      opCodes[613] <= 162;
      opCodes[776] <= 162;
      opCodes[814] <= 162;
      opCodes[852] <= 162;
      opCodes[890] <= 162;
      opCodes[928] <= 162;
      opCodes[970] <= 162;
      opCodes[1008] <= 162;
      opCodes[1046] <= 162;
      opCodes[1084] <= 162;
      opCodes[1122] <= 162;
      opCodes[1501] <= 162;
      opCodes[1539] <= 162;
      opCodes[1577] <= 162;
      opCodes[1615] <= 162;
      opCodes[2017] <= 162;
      opCodes[2058] <= 162;
      opCodes[2099] <= 162;
      opCodes[2140] <= 162;
      opCodes[2181] <= 162;
      opCodes[2222] <= 162;
      opCodes[2263] <= 162;
      opCodes[2304] <= 162;
      opCodes[2345] <= 162;
      opCodes[2386] <= 162;
      opCodes[2427] <= 162;
      opCodes[2468] <= 162;
      opCodes[2509] <= 162;
      opCodes[2550] <= 162;
      opCodes[2591] <= 162;
      opCodes[2632] <= 162;
      opCodes[2772] <= 162;
      opCodes[2813] <= 162;
      opCodes[2854] <= 162;
      opCodes[2895] <= 162;
      opCodes[2936] <= 162;
      opCodes[2977] <= 162;
      opCodes[3018] <= 162;
      opCodes[3059] <= 162;
      opCodes[3100] <= 162;
      opCodes[3165] <= 162;
      opCodes[3206] <= 162;
      opCodes[3247] <= 162;
      opCodes[3288] <= 162;
      opCodes[3329] <= 162;
      opCodes[3370] <= 162;
      opCodes[3411] <= 162;
      opCodes[3452] <= 162;
      opCodes[3493] <= 162;
      opCodes[4646] <= 162;
      opCodes[4687] <= 162;
      opCodes[4728] <= 162;
      opCodes[4769] <= 162;
      opCodes[4810] <= 162;
      opCodes[4851] <= 162;
      opCodes[4892] <= 162;
      opCodes[4933] <= 162;
      opCodes[5045] <= 162;
      opCodes[5086] <= 162;
      opCodes[5127] <= 162;
      opCodes[5168] <= 162;
      opCodes[5209] <= 162;
      opCodes[5250] <= 162;
      opCodes[5291] <= 162;
      opCodes[5332] <= 162;
      opCodes[5373] <= 162;
      opCodes[5606] <= 162;
      opCodes[5644] <= 162;
      opCodes[5682] <= 162;
      opCodes[5720] <= 162;
      opCodes[5758] <= 162;
      opCodes[348] <= 163;
      opCodes[386] <= 163;
      opCodes[424] <= 163;
      opCodes[462] <= 163;
      opCodes[500] <= 163;
      opCodes[538] <= 163;
      opCodes[576] <= 163;
      opCodes[614] <= 163;
      opCodes[777] <= 163;
      opCodes[815] <= 163;
      opCodes[853] <= 163;
      opCodes[891] <= 163;
      opCodes[929] <= 163;
      opCodes[971] <= 163;
      opCodes[1009] <= 163;
      opCodes[1047] <= 163;
      opCodes[1085] <= 163;
      opCodes[1123] <= 163;
      opCodes[1502] <= 163;
      opCodes[1540] <= 163;
      opCodes[1578] <= 163;
      opCodes[1616] <= 163;
      opCodes[2018] <= 163;
      opCodes[2059] <= 163;
      opCodes[2100] <= 163;
      opCodes[2141] <= 163;
      opCodes[2182] <= 163;
      opCodes[2223] <= 163;
      opCodes[2264] <= 163;
      opCodes[2305] <= 163;
      opCodes[2346] <= 163;
      opCodes[2387] <= 163;
      opCodes[2428] <= 163;
      opCodes[2469] <= 163;
      opCodes[2510] <= 163;
      opCodes[2551] <= 163;
      opCodes[2592] <= 163;
      opCodes[2633] <= 163;
      opCodes[2773] <= 163;
      opCodes[2814] <= 163;
      opCodes[2855] <= 163;
      opCodes[2896] <= 163;
      opCodes[2937] <= 163;
      opCodes[2978] <= 163;
      opCodes[3019] <= 163;
      opCodes[3060] <= 163;
      opCodes[3101] <= 163;
      opCodes[3166] <= 163;
      opCodes[3207] <= 163;
      opCodes[3248] <= 163;
      opCodes[3289] <= 163;
      opCodes[3330] <= 163;
      opCodes[3371] <= 163;
      opCodes[3412] <= 163;
      opCodes[3453] <= 163;
      opCodes[3494] <= 163;
      opCodes[4647] <= 163;
      opCodes[4688] <= 163;
      opCodes[4729] <= 163;
      opCodes[4770] <= 163;
      opCodes[4811] <= 163;
      opCodes[4852] <= 163;
      opCodes[4893] <= 163;
      opCodes[4934] <= 163;
      opCodes[5046] <= 163;
      opCodes[5087] <= 163;
      opCodes[5128] <= 163;
      opCodes[5169] <= 163;
      opCodes[5210] <= 163;
      opCodes[5251] <= 163;
      opCodes[5292] <= 163;
      opCodes[5333] <= 163;
      opCodes[5374] <= 163;
      opCodes[5607] <= 163;
      opCodes[5645] <= 163;
      opCodes[5683] <= 163;
      opCodes[5721] <= 163;
      opCodes[5759] <= 163;
      opCodes[349] <= 164;
      opCodes[387] <= 164;
      opCodes[425] <= 164;
      opCodes[463] <= 164;
      opCodes[501] <= 164;
      opCodes[539] <= 164;
      opCodes[577] <= 164;
      opCodes[615] <= 164;
      opCodes[778] <= 164;
      opCodes[816] <= 164;
      opCodes[854] <= 164;
      opCodes[892] <= 164;
      opCodes[930] <= 164;
      opCodes[972] <= 164;
      opCodes[1010] <= 164;
      opCodes[1048] <= 164;
      opCodes[1086] <= 164;
      opCodes[1124] <= 164;
      opCodes[1503] <= 164;
      opCodes[1541] <= 164;
      opCodes[1579] <= 164;
      opCodes[1617] <= 164;
      opCodes[2019] <= 164;
      opCodes[2060] <= 164;
      opCodes[2101] <= 164;
      opCodes[2142] <= 164;
      opCodes[2183] <= 164;
      opCodes[2224] <= 164;
      opCodes[2265] <= 164;
      opCodes[2306] <= 164;
      opCodes[2347] <= 164;
      opCodes[2388] <= 164;
      opCodes[2429] <= 164;
      opCodes[2470] <= 164;
      opCodes[2511] <= 164;
      opCodes[2552] <= 164;
      opCodes[2593] <= 164;
      opCodes[2634] <= 164;
      opCodes[2774] <= 164;
      opCodes[2815] <= 164;
      opCodes[2856] <= 164;
      opCodes[2897] <= 164;
      opCodes[2938] <= 164;
      opCodes[2979] <= 164;
      opCodes[3020] <= 164;
      opCodes[3061] <= 164;
      opCodes[3102] <= 164;
      opCodes[3167] <= 164;
      opCodes[3208] <= 164;
      opCodes[3249] <= 164;
      opCodes[3290] <= 164;
      opCodes[3331] <= 164;
      opCodes[3372] <= 164;
      opCodes[3413] <= 164;
      opCodes[3454] <= 164;
      opCodes[3495] <= 164;
      opCodes[4648] <= 164;
      opCodes[4689] <= 164;
      opCodes[4730] <= 164;
      opCodes[4771] <= 164;
      opCodes[4812] <= 164;
      opCodes[4853] <= 164;
      opCodes[4894] <= 164;
      opCodes[4935] <= 164;
      opCodes[5047] <= 164;
      opCodes[5088] <= 164;
      opCodes[5129] <= 164;
      opCodes[5170] <= 164;
      opCodes[5211] <= 164;
      opCodes[5252] <= 164;
      opCodes[5293] <= 164;
      opCodes[5334] <= 164;
      opCodes[5375] <= 164;
      opCodes[5608] <= 164;
      opCodes[5646] <= 164;
      opCodes[5684] <= 164;
      opCodes[5722] <= 164;
      opCodes[5760] <= 164;
      opCodes[350] <= 165;
      opCodes[388] <= 165;
      opCodes[426] <= 165;
      opCodes[464] <= 165;
      opCodes[502] <= 165;
      opCodes[540] <= 165;
      opCodes[578] <= 165;
      opCodes[616] <= 165;
      opCodes[779] <= 165;
      opCodes[817] <= 165;
      opCodes[855] <= 165;
      opCodes[893] <= 165;
      opCodes[931] <= 165;
      opCodes[973] <= 165;
      opCodes[1011] <= 165;
      opCodes[1049] <= 165;
      opCodes[1087] <= 165;
      opCodes[1125] <= 165;
      opCodes[1504] <= 165;
      opCodes[1542] <= 165;
      opCodes[1580] <= 165;
      opCodes[1618] <= 165;
      opCodes[2020] <= 165;
      opCodes[2061] <= 165;
      opCodes[2102] <= 165;
      opCodes[2143] <= 165;
      opCodes[2184] <= 165;
      opCodes[2225] <= 165;
      opCodes[2266] <= 165;
      opCodes[2307] <= 165;
      opCodes[2348] <= 165;
      opCodes[2389] <= 165;
      opCodes[2430] <= 165;
      opCodes[2471] <= 165;
      opCodes[2512] <= 165;
      opCodes[2553] <= 165;
      opCodes[2594] <= 165;
      opCodes[2635] <= 165;
      opCodes[2775] <= 165;
      opCodes[2816] <= 165;
      opCodes[2857] <= 165;
      opCodes[2898] <= 165;
      opCodes[2939] <= 165;
      opCodes[2980] <= 165;
      opCodes[3021] <= 165;
      opCodes[3062] <= 165;
      opCodes[3103] <= 165;
      opCodes[3168] <= 165;
      opCodes[3209] <= 165;
      opCodes[3250] <= 165;
      opCodes[3291] <= 165;
      opCodes[3332] <= 165;
      opCodes[3373] <= 165;
      opCodes[3414] <= 165;
      opCodes[3455] <= 165;
      opCodes[3496] <= 165;
      opCodes[4649] <= 165;
      opCodes[4690] <= 165;
      opCodes[4731] <= 165;
      opCodes[4772] <= 165;
      opCodes[4813] <= 165;
      opCodes[4854] <= 165;
      opCodes[4895] <= 165;
      opCodes[4936] <= 165;
      opCodes[5048] <= 165;
      opCodes[5089] <= 165;
      opCodes[5130] <= 165;
      opCodes[5171] <= 165;
      opCodes[5212] <= 165;
      opCodes[5253] <= 165;
      opCodes[5294] <= 165;
      opCodes[5335] <= 165;
      opCodes[5376] <= 165;
      opCodes[5609] <= 165;
      opCodes[5647] <= 165;
      opCodes[5685] <= 165;
      opCodes[5723] <= 165;
      opCodes[5761] <= 165;
      opCodes[351] <= 166;
      opCodes[389] <= 166;
      opCodes[427] <= 166;
      opCodes[465] <= 166;
      opCodes[503] <= 166;
      opCodes[541] <= 166;
      opCodes[579] <= 166;
      opCodes[617] <= 166;
      opCodes[780] <= 166;
      opCodes[818] <= 166;
      opCodes[856] <= 166;
      opCodes[894] <= 166;
      opCodes[932] <= 166;
      opCodes[974] <= 166;
      opCodes[1012] <= 166;
      opCodes[1050] <= 166;
      opCodes[1088] <= 166;
      opCodes[1126] <= 166;
      opCodes[1505] <= 166;
      opCodes[1543] <= 166;
      opCodes[1581] <= 166;
      opCodes[1619] <= 166;
      opCodes[2021] <= 166;
      opCodes[2062] <= 166;
      opCodes[2103] <= 166;
      opCodes[2144] <= 166;
      opCodes[2185] <= 166;
      opCodes[2226] <= 166;
      opCodes[2267] <= 166;
      opCodes[2308] <= 166;
      opCodes[2349] <= 166;
      opCodes[2390] <= 166;
      opCodes[2431] <= 166;
      opCodes[2472] <= 166;
      opCodes[2513] <= 166;
      opCodes[2554] <= 166;
      opCodes[2595] <= 166;
      opCodes[2636] <= 166;
      opCodes[2776] <= 166;
      opCodes[2817] <= 166;
      opCodes[2858] <= 166;
      opCodes[2899] <= 166;
      opCodes[2940] <= 166;
      opCodes[2981] <= 166;
      opCodes[3022] <= 166;
      opCodes[3063] <= 166;
      opCodes[3104] <= 166;
      opCodes[3169] <= 166;
      opCodes[3210] <= 166;
      opCodes[3251] <= 166;
      opCodes[3292] <= 166;
      opCodes[3333] <= 166;
      opCodes[3374] <= 166;
      opCodes[3415] <= 166;
      opCodes[3456] <= 166;
      opCodes[3497] <= 166;
      opCodes[4650] <= 166;
      opCodes[4691] <= 166;
      opCodes[4732] <= 166;
      opCodes[4773] <= 166;
      opCodes[4814] <= 166;
      opCodes[4855] <= 166;
      opCodes[4896] <= 166;
      opCodes[4937] <= 166;
      opCodes[5049] <= 166;
      opCodes[5090] <= 166;
      opCodes[5131] <= 166;
      opCodes[5172] <= 166;
      opCodes[5213] <= 166;
      opCodes[5254] <= 166;
      opCodes[5295] <= 166;
      opCodes[5336] <= 166;
      opCodes[5377] <= 166;
      opCodes[5610] <= 166;
      opCodes[5648] <= 166;
      opCodes[5686] <= 166;
      opCodes[5724] <= 166;
      opCodes[5762] <= 166;
      opCodes[353] <= 167;
      opCodes[391] <= 167;
      opCodes[429] <= 167;
      opCodes[467] <= 167;
      opCodes[505] <= 167;
      opCodes[543] <= 167;
      opCodes[581] <= 167;
      opCodes[619] <= 167;
      opCodes[782] <= 167;
      opCodes[820] <= 167;
      opCodes[858] <= 167;
      opCodes[896] <= 167;
      opCodes[934] <= 167;
      opCodes[976] <= 167;
      opCodes[1014] <= 167;
      opCodes[1052] <= 167;
      opCodes[1090] <= 167;
      opCodes[1128] <= 167;
      opCodes[1507] <= 167;
      opCodes[1545] <= 167;
      opCodes[1583] <= 167;
      opCodes[1621] <= 167;
      opCodes[2023] <= 167;
      opCodes[2064] <= 167;
      opCodes[2105] <= 167;
      opCodes[2146] <= 167;
      opCodes[2187] <= 167;
      opCodes[2228] <= 167;
      opCodes[2269] <= 167;
      opCodes[2310] <= 167;
      opCodes[2351] <= 167;
      opCodes[2392] <= 167;
      opCodes[2433] <= 167;
      opCodes[2474] <= 167;
      opCodes[2515] <= 167;
      opCodes[2556] <= 167;
      opCodes[2597] <= 167;
      opCodes[2638] <= 167;
      opCodes[2778] <= 167;
      opCodes[2819] <= 167;
      opCodes[2860] <= 167;
      opCodes[2901] <= 167;
      opCodes[2942] <= 167;
      opCodes[2983] <= 167;
      opCodes[3024] <= 167;
      opCodes[3065] <= 167;
      opCodes[3106] <= 167;
      opCodes[3171] <= 167;
      opCodes[3212] <= 167;
      opCodes[3253] <= 167;
      opCodes[3294] <= 167;
      opCodes[3335] <= 167;
      opCodes[3376] <= 167;
      opCodes[3417] <= 167;
      opCodes[3458] <= 167;
      opCodes[3499] <= 167;
      opCodes[4652] <= 167;
      opCodes[4693] <= 167;
      opCodes[4734] <= 167;
      opCodes[4775] <= 167;
      opCodes[4816] <= 167;
      opCodes[4857] <= 167;
      opCodes[4898] <= 167;
      opCodes[4939] <= 167;
      opCodes[5051] <= 167;
      opCodes[5092] <= 167;
      opCodes[5133] <= 167;
      opCodes[5174] <= 167;
      opCodes[5215] <= 167;
      opCodes[5256] <= 167;
      opCodes[5297] <= 167;
      opCodes[5338] <= 167;
      opCodes[5379] <= 167;
      opCodes[5612] <= 167;
      opCodes[5650] <= 167;
      opCodes[5688] <= 167;
      opCodes[5726] <= 167;
      opCodes[5764] <= 167;
      opCodes[354] <= 168;
      opCodes[392] <= 168;
      opCodes[430] <= 168;
      opCodes[468] <= 168;
      opCodes[506] <= 168;
      opCodes[544] <= 168;
      opCodes[582] <= 168;
      opCodes[620] <= 168;
      opCodes[783] <= 168;
      opCodes[821] <= 168;
      opCodes[859] <= 168;
      opCodes[897] <= 168;
      opCodes[935] <= 168;
      opCodes[977] <= 168;
      opCodes[1015] <= 168;
      opCodes[1053] <= 168;
      opCodes[1091] <= 168;
      opCodes[1129] <= 168;
      opCodes[1508] <= 168;
      opCodes[1546] <= 168;
      opCodes[1584] <= 168;
      opCodes[1622] <= 168;
      opCodes[2024] <= 168;
      opCodes[2065] <= 168;
      opCodes[2106] <= 168;
      opCodes[2147] <= 168;
      opCodes[2188] <= 168;
      opCodes[2229] <= 168;
      opCodes[2270] <= 168;
      opCodes[2311] <= 168;
      opCodes[2352] <= 168;
      opCodes[2393] <= 168;
      opCodes[2434] <= 168;
      opCodes[2475] <= 168;
      opCodes[2516] <= 168;
      opCodes[2557] <= 168;
      opCodes[2598] <= 168;
      opCodes[2639] <= 168;
      opCodes[2779] <= 168;
      opCodes[2820] <= 168;
      opCodes[2861] <= 168;
      opCodes[2902] <= 168;
      opCodes[2943] <= 168;
      opCodes[2984] <= 168;
      opCodes[3025] <= 168;
      opCodes[3066] <= 168;
      opCodes[3107] <= 168;
      opCodes[3172] <= 168;
      opCodes[3213] <= 168;
      opCodes[3254] <= 168;
      opCodes[3295] <= 168;
      opCodes[3336] <= 168;
      opCodes[3377] <= 168;
      opCodes[3418] <= 168;
      opCodes[3459] <= 168;
      opCodes[3500] <= 168;
      opCodes[4653] <= 168;
      opCodes[4694] <= 168;
      opCodes[4735] <= 168;
      opCodes[4776] <= 168;
      opCodes[4817] <= 168;
      opCodes[4858] <= 168;
      opCodes[4899] <= 168;
      opCodes[4940] <= 168;
      opCodes[5052] <= 168;
      opCodes[5093] <= 168;
      opCodes[5134] <= 168;
      opCodes[5175] <= 168;
      opCodes[5216] <= 168;
      opCodes[5257] <= 168;
      opCodes[5298] <= 168;
      opCodes[5339] <= 168;
      opCodes[5380] <= 168;
      opCodes[5613] <= 168;
      opCodes[5651] <= 168;
      opCodes[5689] <= 168;
      opCodes[5727] <= 168;
      opCodes[5765] <= 168;
      opCodes[356] <= 169;
      opCodes[394] <= 169;
      opCodes[432] <= 169;
      opCodes[470] <= 169;
      opCodes[508] <= 169;
      opCodes[546] <= 169;
      opCodes[584] <= 169;
      opCodes[622] <= 169;
      opCodes[785] <= 169;
      opCodes[823] <= 169;
      opCodes[861] <= 169;
      opCodes[899] <= 169;
      opCodes[937] <= 169;
      opCodes[979] <= 169;
      opCodes[1017] <= 169;
      opCodes[1055] <= 169;
      opCodes[1093] <= 169;
      opCodes[1131] <= 169;
      opCodes[1510] <= 169;
      opCodes[1548] <= 169;
      opCodes[1586] <= 169;
      opCodes[1624] <= 169;
      opCodes[2026] <= 169;
      opCodes[2067] <= 169;
      opCodes[2108] <= 169;
      opCodes[2149] <= 169;
      opCodes[2190] <= 169;
      opCodes[2231] <= 169;
      opCodes[2272] <= 169;
      opCodes[2313] <= 169;
      opCodes[2354] <= 169;
      opCodes[2395] <= 169;
      opCodes[2436] <= 169;
      opCodes[2477] <= 169;
      opCodes[2518] <= 169;
      opCodes[2559] <= 169;
      opCodes[2600] <= 169;
      opCodes[2641] <= 169;
      opCodes[2781] <= 169;
      opCodes[2822] <= 169;
      opCodes[2863] <= 169;
      opCodes[2904] <= 169;
      opCodes[2945] <= 169;
      opCodes[2986] <= 169;
      opCodes[3027] <= 169;
      opCodes[3068] <= 169;
      opCodes[3109] <= 169;
      opCodes[3174] <= 169;
      opCodes[3215] <= 169;
      opCodes[3256] <= 169;
      opCodes[3297] <= 169;
      opCodes[3338] <= 169;
      opCodes[3379] <= 169;
      opCodes[3420] <= 169;
      opCodes[3461] <= 169;
      opCodes[3502] <= 169;
      opCodes[4655] <= 169;
      opCodes[4696] <= 169;
      opCodes[4737] <= 169;
      opCodes[4778] <= 169;
      opCodes[4819] <= 169;
      opCodes[4860] <= 169;
      opCodes[4901] <= 169;
      opCodes[4942] <= 169;
      opCodes[5054] <= 169;
      opCodes[5095] <= 169;
      opCodes[5136] <= 169;
      opCodes[5177] <= 169;
      opCodes[5218] <= 169;
      opCodes[5259] <= 169;
      opCodes[5300] <= 169;
      opCodes[5341] <= 169;
      opCodes[5382] <= 169;
      opCodes[5615] <= 169;
      opCodes[5653] <= 169;
      opCodes[5691] <= 169;
      opCodes[5729] <= 169;
      opCodes[5767] <= 169;
      opCodes[357] <= 170;
      opCodes[384] <= 171;
      opCodes[395] <= 172;
      opCodes[422] <= 173;
      opCodes[433] <= 174;
      opCodes[460] <= 175;
      opCodes[471] <= 176;
      opCodes[498] <= 177;
      opCodes[509] <= 178;
      opCodes[536] <= 179;
      opCodes[547] <= 180;
      opCodes[574] <= 181;
      opCodes[585] <= 182;
      opCodes[612] <= 183;
      opCodes[623] <= 184;
      opCodes[644] <= 185;
      opCodes[657] <= 186;
      opCodes[658] <= 187;
      opCodes[659] <= 188;
      opCodes[661] <= 188;
      opCodes[664] <= 188;
      opCodes[660] <= 189;
      opCodes[662] <= 190;
      opCodes[669] <= 190;
      opCodes[663] <= 191;
      opCodes[1667] <= 191;
      opCodes[665] <= 192;
      opCodes[668] <= 193;
      opCodes[1151] <= 193;
      opCodes[2000] <= 193;
      opCodes[2755] <= 193;
      opCodes[696] <= 194;
      opCodes[698] <= 195;
      opCodes[699] <= 196;
      opCodes[727] <= 196;
      opCodes[790] <= 196;
      opCodes[828] <= 196;
      opCodes[866] <= 196;
      opCodes[904] <= 196;
      opCodes[944] <= 196;
      opCodes[1154] <= 196;
      opCodes[700] <= 197;
      opCodes[702] <= 198;
      opCodes[704] <= 199;
      opCodes[705] <= 200;
      opCodes[706] <= 201;
      opCodes[728] <= 202;
      opCodes[761] <= 202;
      opCodes[5591] <= 202;
      opCodes[729] <= 203;
      opCodes[762] <= 203;
      opCodes[5592] <= 203;
      opCodes[731] <= 204;
      opCodes[732] <= 205;
      opCodes[760] <= 205;
      opCodes[984] <= 205;
      opCodes[1022] <= 205;
      opCodes[1060] <= 205;
      opCodes[1098] <= 205;
      opCodes[1136] <= 205;
      opCodes[1167] <= 205;
      opCodes[733] <= 206;
      opCodes[735] <= 207;
      opCodes[737] <= 208;
      opCodes[738] <= 209;
      opCodes[739] <= 210;
      opCodes[775] <= 211;
      opCodes[786] <= 212;
      opCodes[813] <= 213;
      opCodes[824] <= 214;
      opCodes[851] <= 215;
      opCodes[862] <= 216;
      opCodes[889] <= 217;
      opCodes[900] <= 218;
      opCodes[927] <= 219;
      opCodes[938] <= 220;
      opCodes[943] <= 221;
      opCodes[969] <= 222;
      opCodes[980] <= 223;
      opCodes[1007] <= 224;
      opCodes[1018] <= 225;
      opCodes[1045] <= 226;
      opCodes[1056] <= 227;
      opCodes[1083] <= 228;
      opCodes[1094] <= 229;
      opCodes[1121] <= 230;
      opCodes[1132] <= 231;
      opCodes[1152] <= 232;
      opCodes[1183] <= 233;
      opCodes[1192] <= 234;
      opCodes[1205] <= 234;
      opCodes[1194] <= 235;
      opCodes[1200] <= 236;
      opCodes[1206] <= 237;
      opCodes[1217] <= 238;
      opCodes[1296] <= 238;
      opCodes[1233] <= 239;
      opCodes[1246] <= 239;
      opCodes[1235] <= 240;
      opCodes[1241] <= 241;
      opCodes[1247] <= 242;
      opCodes[1259] <= 243;
      opCodes[1269] <= 244;
      opCodes[1282] <= 244;
      opCodes[1271] <= 245;
      opCodes[1277] <= 246;
      opCodes[1283] <= 247;
      opCodes[1304] <= 248;
      opCodes[1305] <= 249;
      opCodes[1308] <= 250;
      opCodes[1322] <= 251;
      opCodes[1328] <= 252;
      opCodes[1402] <= 252;
      opCodes[1340] <= 253;
      opCodes[1350] <= 254;
      opCodes[1363] <= 254;
      opCodes[1352] <= 255;
      opCodes[1358] <= 256;
      opCodes[1364] <= 257;
      opCodes[1381] <= 258;
      opCodes[1392] <= 259;
      opCodes[1409] <= 260;
      opCodes[1422] <= 261;
      opCodes[1435] <= 261;
      opCodes[1424] <= 262;
      opCodes[1430] <= 263;
      opCodes[1436] <= 264;
      opCodes[1448] <= 265;
      opCodes[1450] <= 266;
      opCodes[1452] <= 267;
      opCodes[1454] <= 268;
      opCodes[1456] <= 269;
      opCodes[1457] <= 270;
      opCodes[1485] <= 270;
      opCodes[1515] <= 270;
      opCodes[1553] <= 270;
      opCodes[1591] <= 270;
      opCodes[1629] <= 270;
      opCodes[1649] <= 270;
      opCodes[1673] <= 270;
      opCodes[1458] <= 271;
      opCodes[1460] <= 272;
      opCodes[1462] <= 273;
      opCodes[1463] <= 274;
      opCodes[1464] <= 275;
      opCodes[1488] <= 276;
      opCodes[1526] <= 276;
      opCodes[1564] <= 276;
      opCodes[1602] <= 276;
      opCodes[1640] <= 276;
      opCodes[1500] <= 277;
      opCodes[1511] <= 278;
      opCodes[1538] <= 279;
      opCodes[1549] <= 280;
      opCodes[1576] <= 281;
      opCodes[1587] <= 282;
      opCodes[1614] <= 283;
      opCodes[1625] <= 284;
      opCodes[1648] <= 285;
      opCodes[1661] <= 286;
      opCodes[1662] <= 287;
      opCodes[1663] <= 288;
      opCodes[1665] <= 288;
      opCodes[1668] <= 288;
      opCodes[1664] <= 289;
      opCodes[1666] <= 290;
      opCodes[1671] <= 290;
      opCodes[1669] <= 291;
      opCodes[1675] <= 292;
      opCodes[1687] <= 293;
      opCodes[1698] <= 294;
      opCodes[1711] <= 295;
      opCodes[1720] <= 296;
      opCodes[1733] <= 296;
      opCodes[1722] <= 297;
      opCodes[1728] <= 298;
      opCodes[1734] <= 299;
      opCodes[1745] <= 300;
      opCodes[1824] <= 300;
      opCodes[1761] <= 301;
      opCodes[1774] <= 301;
      opCodes[1763] <= 302;
      opCodes[1769] <= 303;
      opCodes[1775] <= 304;
      opCodes[1787] <= 305;
      opCodes[1797] <= 306;
      opCodes[1810] <= 306;
      opCodes[1799] <= 307;
      opCodes[1805] <= 308;
      opCodes[1811] <= 309;
      opCodes[1832] <= 310;
      opCodes[1833] <= 311;
      opCodes[1836] <= 312;
      opCodes[1850] <= 313;
      opCodes[1856] <= 314;
      opCodes[1930] <= 314;
      opCodes[1868] <= 315;
      opCodes[1878] <= 316;
      opCodes[1891] <= 316;
      opCodes[1880] <= 317;
      opCodes[1886] <= 318;
      opCodes[1892] <= 319;
      opCodes[1909] <= 320;
      opCodes[1920] <= 321;
      opCodes[1934] <= 322;
      opCodes[1938] <= 323;
      opCodes[1949] <= 323;
      opCodes[1997] <= 323;
      opCodes[2717] <= 323;
      opCodes[2745] <= 323;
      opCodes[1939] <= 324;
      opCodes[1946] <= 325;
      opCodes[1947] <= 326;
      opCodes[1948] <= 327;
      opCodes[2043] <= 327;
      opCodes[2371] <= 327;
      opCodes[2798] <= 327;
      opCodes[3191] <= 327;
      opCodes[3735] <= 327;
      opCodes[4169] <= 327;
      opCodes[4672] <= 327;
      opCodes[5071] <= 327;
      opCodes[1957] <= 328;
      opCodes[1968] <= 329;
      opCodes[1970] <= 330;
      opCodes[1976] <= 330;
      opCodes[3663] <= 330;
      opCodes[3669] <= 330;
      opCodes[4600] <= 330;
      opCodes[4606] <= 330;
      opCodes[1971] <= 331;
      opCodes[3664] <= 331;
      opCodes[4601] <= 331;
      opCodes[1977] <= 332;
      opCodes[2716] <= 332;
      opCodes[3670] <= 332;
      opCodes[4021] <= 332;
      opCodes[4607] <= 332;
      opCodes[4958] <= 332;
      opCodes[1978] <= 333;
      opCodes[1979] <= 334;
      opCodes[2004] <= 334;
      opCodes[2045] <= 334;
      opCodes[2086] <= 334;
      opCodes[2127] <= 334;
      opCodes[2168] <= 334;
      opCodes[2209] <= 334;
      opCodes[2250] <= 334;
      opCodes[2291] <= 334;
      opCodes[2660] <= 334;
      opCodes[2686] <= 334;
      opCodes[2718] <= 334;
      opCodes[2759] <= 334;
      opCodes[2800] <= 334;
      opCodes[2841] <= 334;
      opCodes[2882] <= 334;
      opCodes[2923] <= 334;
      opCodes[2964] <= 334;
      opCodes[3005] <= 334;
      opCodes[3046] <= 334;
      opCodes[3087] <= 334;
      opCodes[3125] <= 334;
      opCodes[3542] <= 334;
      opCodes[3568] <= 334;
      opCodes[1984] <= 335;
      opCodes[2726] <= 335;
      opCodes[1985] <= 336;
      opCodes[2332] <= 336;
      opCodes[2373] <= 336;
      opCodes[2414] <= 336;
      opCodes[2455] <= 336;
      opCodes[2496] <= 336;
      opCodes[2537] <= 336;
      opCodes[2578] <= 336;
      opCodes[2619] <= 336;
      opCodes[2688] <= 336;
      opCodes[2714] <= 336;
      opCodes[2727] <= 336;
      opCodes[3152] <= 336;
      opCodes[3193] <= 336;
      opCodes[3234] <= 336;
      opCodes[3275] <= 336;
      opCodes[3316] <= 336;
      opCodes[3357] <= 336;
      opCodes[3398] <= 336;
      opCodes[3439] <= 336;
      opCodes[3480] <= 336;
      opCodes[3518] <= 336;
      opCodes[3570] <= 336;
      opCodes[3596] <= 336;
      opCodes[1990] <= 337;
      opCodes[2735] <= 337;
      opCodes[1991] <= 338;
      opCodes[2001] <= 338;
      opCodes[2042] <= 338;
      opCodes[2083] <= 338;
      opCodes[2124] <= 338;
      opCodes[2165] <= 338;
      opCodes[2206] <= 338;
      opCodes[2247] <= 338;
      opCodes[2288] <= 338;
      opCodes[2736] <= 338;
      opCodes[2756] <= 338;
      opCodes[2797] <= 338;
      opCodes[2838] <= 338;
      opCodes[2879] <= 338;
      opCodes[2920] <= 338;
      opCodes[2961] <= 338;
      opCodes[3002] <= 338;
      opCodes[3043] <= 338;
      opCodes[3084] <= 338;
      opCodes[1992] <= 339;
      opCodes[1994] <= 339;
      opCodes[2737] <= 339;
      opCodes[2739] <= 339;
      opCodes[2742] <= 339;
      opCodes[1993] <= 340;
      opCodes[2738] <= 340;
      opCodes[1995] <= 341;
      opCodes[2740] <= 341;
      opCodes[2743] <= 341;
      opCodes[2002] <= 342;
      opCodes[2330] <= 342;
      opCodes[2757] <= 342;
      opCodes[3150] <= 342;
      opCodes[3694] <= 342;
      opCodes[4128] <= 342;
      opCodes[4631] <= 342;
      opCodes[5030] <= 342;
      opCodes[2003] <= 343;
      opCodes[2044] <= 343;
      opCodes[2085] <= 343;
      opCodes[2126] <= 343;
      opCodes[2167] <= 343;
      opCodes[2208] <= 343;
      opCodes[2249] <= 343;
      opCodes[2290] <= 343;
      opCodes[2016] <= 344;
      opCodes[2027] <= 345;
      opCodes[2057] <= 346;
      opCodes[2068] <= 347;
      opCodes[2084] <= 348;
      opCodes[2412] <= 348;
      opCodes[2839] <= 348;
      opCodes[3232] <= 348;
      opCodes[3776] <= 348;
      opCodes[4210] <= 348;
      opCodes[4713] <= 348;
      opCodes[5112] <= 348;
      opCodes[2098] <= 349;
      opCodes[2109] <= 350;
      opCodes[2125] <= 351;
      opCodes[2453] <= 351;
      opCodes[2880] <= 351;
      opCodes[3273] <= 351;
      opCodes[3817] <= 351;
      opCodes[4251] <= 351;
      opCodes[4754] <= 351;
      opCodes[5153] <= 351;
      opCodes[2139] <= 352;
      opCodes[2150] <= 353;
      opCodes[2166] <= 354;
      opCodes[2494] <= 354;
      opCodes[2921] <= 354;
      opCodes[3314] <= 354;
      opCodes[3858] <= 354;
      opCodes[4292] <= 354;
      opCodes[4795] <= 354;
      opCodes[5194] <= 354;
      opCodes[2180] <= 355;
      opCodes[2191] <= 356;
      opCodes[2207] <= 357;
      opCodes[2535] <= 357;
      opCodes[2962] <= 357;
      opCodes[3355] <= 357;
      opCodes[3899] <= 357;
      opCodes[4333] <= 357;
      opCodes[4836] <= 357;
      opCodes[5235] <= 357;
      opCodes[2221] <= 358;
      opCodes[2232] <= 359;
      opCodes[2248] <= 360;
      opCodes[2576] <= 360;
      opCodes[3003] <= 360;
      opCodes[3396] <= 360;
      opCodes[3940] <= 360;
      opCodes[4374] <= 360;
      opCodes[4877] <= 360;
      opCodes[5276] <= 360;
      opCodes[2262] <= 361;
      opCodes[2273] <= 362;
      opCodes[2289] <= 363;
      opCodes[2617] <= 363;
      opCodes[3044] <= 363;
      opCodes[3437] <= 363;
      opCodes[3981] <= 363;
      opCodes[4415] <= 363;
      opCodes[4918] <= 363;
      opCodes[5317] <= 363;
      opCodes[2303] <= 364;
      opCodes[2314] <= 365;
      opCodes[2329] <= 366;
      opCodes[2370] <= 366;
      opCodes[2411] <= 366;
      opCodes[2452] <= 366;
      opCodes[2493] <= 366;
      opCodes[2534] <= 366;
      opCodes[2575] <= 366;
      opCodes[2616] <= 366;
      opCodes[3149] <= 366;
      opCodes[3190] <= 366;
      opCodes[3231] <= 366;
      opCodes[3272] <= 366;
      opCodes[3313] <= 366;
      opCodes[3354] <= 366;
      opCodes[3395] <= 366;
      opCodes[3436] <= 366;
      opCodes[3477] <= 366;
      opCodes[2331] <= 367;
      opCodes[2372] <= 367;
      opCodes[2413] <= 367;
      opCodes[2454] <= 367;
      opCodes[2495] <= 367;
      opCodes[2536] <= 367;
      opCodes[2577] <= 367;
      opCodes[2618] <= 367;
      opCodes[2344] <= 368;
      opCodes[2355] <= 369;
      opCodes[2385] <= 370;
      opCodes[2396] <= 371;
      opCodes[2426] <= 372;
      opCodes[2437] <= 373;
      opCodes[2467] <= 374;
      opCodes[2478] <= 375;
      opCodes[2508] <= 376;
      opCodes[2519] <= 377;
      opCodes[2549] <= 378;
      opCodes[2560] <= 379;
      opCodes[2590] <= 380;
      opCodes[2601] <= 381;
      opCodes[2631] <= 382;
      opCodes[2642] <= 383;
      opCodes[2661] <= 384;
      opCodes[3543] <= 384;
      opCodes[2662] <= 385;
      opCodes[3544] <= 385;
      opCodes[2663] <= 386;
      opCodes[3545] <= 386;
      opCodes[2664] <= 387;
      opCodes[2692] <= 387;
      opCodes[3546] <= 387;
      opCodes[3574] <= 387;
      opCodes[4500] <= 387;
      opCodes[5402] <= 387;
      opCodes[2665] <= 388;
      opCodes[2693] <= 388;
      opCodes[3547] <= 388;
      opCodes[3575] <= 388;
      opCodes[4501] <= 388;
      opCodes[5403] <= 388;
      opCodes[2666] <= 389;
      opCodes[2694] <= 389;
      opCodes[3548] <= 389;
      opCodes[3576] <= 389;
      opCodes[4502] <= 389;
      opCodes[5404] <= 389;
      opCodes[2667] <= 390;
      opCodes[2695] <= 390;
      opCodes[3549] <= 390;
      opCodes[3577] <= 390;
      opCodes[4503] <= 390;
      opCodes[5405] <= 390;
      opCodes[2668] <= 391;
      opCodes[2696] <= 391;
      opCodes[3550] <= 391;
      opCodes[3578] <= 391;
      opCodes[4504] <= 391;
      opCodes[5406] <= 391;
      opCodes[2669] <= 392;
      opCodes[2697] <= 392;
      opCodes[3551] <= 392;
      opCodes[3579] <= 392;
      opCodes[4505] <= 392;
      opCodes[5407] <= 392;
      opCodes[2670] <= 393;
      opCodes[2698] <= 393;
      opCodes[3552] <= 393;
      opCodes[3580] <= 393;
      opCodes[4506] <= 393;
      opCodes[5408] <= 393;
      opCodes[2671] <= 394;
      opCodes[2699] <= 394;
      opCodes[3553] <= 394;
      opCodes[3581] <= 394;
      opCodes[4507] <= 394;
      opCodes[5409] <= 394;
      opCodes[2672] <= 395;
      opCodes[2700] <= 395;
      opCodes[3554] <= 395;
      opCodes[3582] <= 395;
      opCodes[4508] <= 395;
      opCodes[5410] <= 395;
      opCodes[2673] <= 396;
      opCodes[2701] <= 396;
      opCodes[3555] <= 396;
      opCodes[3583] <= 396;
      opCodes[4509] <= 396;
      opCodes[5411] <= 396;
      opCodes[2674] <= 397;
      opCodes[2702] <= 397;
      opCodes[3556] <= 397;
      opCodes[3584] <= 397;
      opCodes[4510] <= 397;
      opCodes[5412] <= 397;
      opCodes[2675] <= 398;
      opCodes[2703] <= 398;
      opCodes[3557] <= 398;
      opCodes[3585] <= 398;
      opCodes[4511] <= 398;
      opCodes[5413] <= 398;
      opCodes[2676] <= 399;
      opCodes[2704] <= 399;
      opCodes[3558] <= 399;
      opCodes[3586] <= 399;
      opCodes[4512] <= 399;
      opCodes[5414] <= 399;
      opCodes[2677] <= 400;
      opCodes[2705] <= 400;
      opCodes[3559] <= 400;
      opCodes[3587] <= 400;
      opCodes[4513] <= 400;
      opCodes[5415] <= 400;
      opCodes[2678] <= 401;
      opCodes[2706] <= 401;
      opCodes[3560] <= 401;
      opCodes[3588] <= 401;
      opCodes[4514] <= 401;
      opCodes[5416] <= 401;
      opCodes[2679] <= 402;
      opCodes[2707] <= 402;
      opCodes[3561] <= 402;
      opCodes[3589] <= 402;
      opCodes[4515] <= 402;
      opCodes[5417] <= 402;
      opCodes[2680] <= 403;
      opCodes[2708] <= 403;
      opCodes[3562] <= 403;
      opCodes[3590] <= 403;
      opCodes[4516] <= 403;
      opCodes[5418] <= 403;
      opCodes[2681] <= 404;
      opCodes[2709] <= 404;
      opCodes[3563] <= 404;
      opCodes[3591] <= 404;
      opCodes[4517] <= 404;
      opCodes[5419] <= 404;
      opCodes[2682] <= 405;
      opCodes[2710] <= 405;
      opCodes[3564] <= 405;
      opCodes[3592] <= 405;
      opCodes[4518] <= 405;
      opCodes[5420] <= 405;
      opCodes[2683] <= 406;
      opCodes[2711] <= 406;
      opCodes[3565] <= 406;
      opCodes[3593] <= 406;
      opCodes[4519] <= 406;
      opCodes[5421] <= 406;
      opCodes[2685] <= 407;
      opCodes[3567] <= 407;
      opCodes[2689] <= 408;
      opCodes[3571] <= 408;
      opCodes[2690] <= 409;
      opCodes[3572] <= 409;
      opCodes[2691] <= 410;
      opCodes[3573] <= 410;
      opCodes[2713] <= 411;
      opCodes[3595] <= 411;
      opCodes[2754] <= 412;
      opCodes[2758] <= 413;
      opCodes[2799] <= 413;
      opCodes[2840] <= 413;
      opCodes[2881] <= 413;
      opCodes[2922] <= 413;
      opCodes[2963] <= 413;
      opCodes[3004] <= 413;
      opCodes[3045] <= 413;
      opCodes[3086] <= 413;
      opCodes[2771] <= 414;
      opCodes[2782] <= 415;
      opCodes[2812] <= 416;
      opCodes[2823] <= 417;
      opCodes[2853] <= 418;
      opCodes[2864] <= 419;
      opCodes[2894] <= 420;
      opCodes[2905] <= 421;
      opCodes[2935] <= 422;
      opCodes[2946] <= 423;
      opCodes[2976] <= 424;
      opCodes[2987] <= 425;
      opCodes[3017] <= 426;
      opCodes[3028] <= 427;
      opCodes[3058] <= 428;
      opCodes[3069] <= 429;
      opCodes[3099] <= 430;
      opCodes[3110] <= 431;
      opCodes[3138] <= 432;
      opCodes[3151] <= 433;
      opCodes[3192] <= 433;
      opCodes[3233] <= 433;
      opCodes[3274] <= 433;
      opCodes[3315] <= 433;
      opCodes[3356] <= 433;
      opCodes[3397] <= 433;
      opCodes[3438] <= 433;
      opCodes[3479] <= 433;
      opCodes[3164] <= 434;
      opCodes[3175] <= 435;
      opCodes[3205] <= 436;
      opCodes[3216] <= 437;
      opCodes[3246] <= 438;
      opCodes[3257] <= 439;
      opCodes[3287] <= 440;
      opCodes[3298] <= 441;
      opCodes[3328] <= 442;
      opCodes[3339] <= 443;
      opCodes[3369] <= 444;
      opCodes[3380] <= 445;
      opCodes[3410] <= 446;
      opCodes[3421] <= 447;
      opCodes[3451] <= 448;
      opCodes[3462] <= 449;
      opCodes[3492] <= 450;
      opCodes[3503] <= 451;
      opCodes[3600] <= 452;
      opCodes[3601] <= 453;
      opCodes[3607] <= 454;
      opCodes[3616] <= 455;
      opCodes[3619] <= 455;
      opCodes[3617] <= 456;
      opCodes[3620] <= 457;
      opCodes[3621] <= 458;
      opCodes[3622] <= 459;
      opCodes[3624] <= 460;
      opCodes[3625] <= 461;
      opCodes[4563] <= 461;
      opCodes[4568] <= 461;
      opCodes[5493] <= 461;
      opCodes[3626] <= 462;
      opCodes[3627] <= 463;
      opCodes[3628] <= 464;
      opCodes[3643] <= 464;
      opCodes[3654] <= 464;
      opCodes[4053] <= 464;
      opCodes[4526] <= 464;
      opCodes[3629] <= 465;
      opCodes[3630] <= 466;
      opCodes[3641] <= 466;
      opCodes[3662] <= 466;
      opCodes[4051] <= 466;
      opCodes[4524] <= 466;
      opCodes[3638] <= 467;
      opCodes[3639] <= 468;
      opCodes[3640] <= 469;
      opCodes[3690] <= 469;
      opCodes[3653] <= 470;
      opCodes[3661] <= 471;
      opCodes[3671] <= 472;
      opCodes[3672] <= 473;
      opCodes[3696] <= 473;
      opCodes[3737] <= 473;
      opCodes[3778] <= 473;
      opCodes[3819] <= 473;
      opCodes[3860] <= 473;
      opCodes[3901] <= 473;
      opCodes[3942] <= 473;
      opCodes[3983] <= 473;
      opCodes[4023] <= 473;
      opCodes[4064] <= 473;
      opCodes[4104] <= 473;
      opCodes[4115] <= 473;
      opCodes[4130] <= 473;
      opCodes[4171] <= 473;
      opCodes[4212] <= 473;
      opCodes[4253] <= 473;
      opCodes[4294] <= 473;
      opCodes[4335] <= 473;
      opCodes[4376] <= 473;
      opCodes[4417] <= 473;
      opCodes[4458] <= 473;
      opCodes[4496] <= 473;
      opCodes[4522] <= 473;
      opCodes[3677] <= 474;
      opCodes[4031] <= 474;
      opCodes[3678] <= 475;
      opCodes[3707] <= 475;
      opCodes[3748] <= 475;
      opCodes[3789] <= 475;
      opCodes[3830] <= 475;
      opCodes[3871] <= 475;
      opCodes[3912] <= 475;
      opCodes[3953] <= 475;
      opCodes[3994] <= 475;
      opCodes[4032] <= 475;
      opCodes[4075] <= 475;
      opCodes[4141] <= 475;
      opCodes[4182] <= 475;
      opCodes[4223] <= 475;
      opCodes[4264] <= 475;
      opCodes[4305] <= 475;
      opCodes[4346] <= 475;
      opCodes[4387] <= 475;
      opCodes[4428] <= 475;
      opCodes[4469] <= 475;
      opCodes[3683] <= 476;
      opCodes[4040] <= 476;
      opCodes[3684] <= 477;
      opCodes[4041] <= 477;
      opCodes[3685] <= 478;
      opCodes[3687] <= 478;
      opCodes[4042] <= 478;
      opCodes[4045] <= 478;
      opCodes[4047] <= 478;
      opCodes[3686] <= 479;
      opCodes[4046] <= 479;
      opCodes[3688] <= 480;
      opCodes[4043] <= 480;
      opCodes[4048] <= 480;
      opCodes[3691] <= 481;
      opCodes[3692] <= 482;
      opCodes[4123] <= 482;
      opCodes[4126] <= 482;
      opCodes[3693] <= 483;
      opCodes[3734] <= 483;
      opCodes[3775] <= 483;
      opCodes[3816] <= 483;
      opCodes[3857] <= 483;
      opCodes[3898] <= 483;
      opCodes[3939] <= 483;
      opCodes[3980] <= 483;
      opCodes[4124] <= 483;
      opCodes[4127] <= 483;
      opCodes[4168] <= 483;
      opCodes[4209] <= 483;
      opCodes[4250] <= 483;
      opCodes[4291] <= 483;
      opCodes[4332] <= 483;
      opCodes[4373] <= 483;
      opCodes[4414] <= 483;
      opCodes[4455] <= 483;
      opCodes[3695] <= 484;
      opCodes[3736] <= 484;
      opCodes[3777] <= 484;
      opCodes[3818] <= 484;
      opCodes[3859] <= 484;
      opCodes[3900] <= 484;
      opCodes[3941] <= 484;
      opCodes[3982] <= 484;
      opCodes[3710] <= 485;
      opCodes[3724] <= 485;
      opCodes[3751] <= 485;
      opCodes[3765] <= 485;
      opCodes[3792] <= 485;
      opCodes[3806] <= 485;
      opCodes[3833] <= 485;
      opCodes[3847] <= 485;
      opCodes[3874] <= 485;
      opCodes[3888] <= 485;
      opCodes[3915] <= 485;
      opCodes[3929] <= 485;
      opCodes[3956] <= 485;
      opCodes[3970] <= 485;
      opCodes[3997] <= 485;
      opCodes[4011] <= 485;
      opCodes[4080] <= 485;
      opCodes[4094] <= 485;
      opCodes[4144] <= 485;
      opCodes[4158] <= 485;
      opCodes[4185] <= 485;
      opCodes[4199] <= 485;
      opCodes[4226] <= 485;
      opCodes[4240] <= 485;
      opCodes[4267] <= 485;
      opCodes[4281] <= 485;
      opCodes[4308] <= 485;
      opCodes[4322] <= 485;
      opCodes[4349] <= 485;
      opCodes[4363] <= 485;
      opCodes[4390] <= 485;
      opCodes[4404] <= 485;
      opCodes[4431] <= 485;
      opCodes[4445] <= 485;
      opCodes[4472] <= 485;
      opCodes[4486] <= 485;
      opCodes[3711] <= 486;
      opCodes[3713] <= 486;
      opCodes[3722] <= 486;
      opCodes[3752] <= 486;
      opCodes[3754] <= 486;
      opCodes[3763] <= 486;
      opCodes[3793] <= 486;
      opCodes[3795] <= 486;
      opCodes[3804] <= 486;
      opCodes[3834] <= 486;
      opCodes[3836] <= 486;
      opCodes[3845] <= 486;
      opCodes[3875] <= 486;
      opCodes[3877] <= 486;
      opCodes[3886] <= 486;
      opCodes[3916] <= 486;
      opCodes[3918] <= 486;
      opCodes[3927] <= 486;
      opCodes[3957] <= 486;
      opCodes[3959] <= 486;
      opCodes[3968] <= 486;
      opCodes[3998] <= 486;
      opCodes[4000] <= 486;
      opCodes[4009] <= 486;
      opCodes[4081] <= 486;
      opCodes[4083] <= 486;
      opCodes[4092] <= 486;
      opCodes[4145] <= 486;
      opCodes[4147] <= 486;
      opCodes[4156] <= 486;
      opCodes[4186] <= 486;
      opCodes[4188] <= 486;
      opCodes[4197] <= 486;
      opCodes[4227] <= 486;
      opCodes[4229] <= 486;
      opCodes[4238] <= 486;
      opCodes[4268] <= 486;
      opCodes[4270] <= 486;
      opCodes[4279] <= 486;
      opCodes[4309] <= 486;
      opCodes[4311] <= 486;
      opCodes[4320] <= 486;
      opCodes[4350] <= 486;
      opCodes[4352] <= 486;
      opCodes[4361] <= 486;
      opCodes[4391] <= 486;
      opCodes[4393] <= 486;
      opCodes[4402] <= 486;
      opCodes[4432] <= 486;
      opCodes[4434] <= 486;
      opCodes[4443] <= 486;
      opCodes[4473] <= 486;
      opCodes[4475] <= 486;
      opCodes[4484] <= 486;
      opCodes[3712] <= 487;
      opCodes[3714] <= 488;
      opCodes[3717] <= 488;
      opCodes[3755] <= 488;
      opCodes[3758] <= 488;
      opCodes[3796] <= 488;
      opCodes[3799] <= 488;
      opCodes[3837] <= 488;
      opCodes[3840] <= 488;
      opCodes[3878] <= 488;
      opCodes[3881] <= 488;
      opCodes[3919] <= 488;
      opCodes[3922] <= 488;
      opCodes[3960] <= 488;
      opCodes[3963] <= 488;
      opCodes[4001] <= 488;
      opCodes[4004] <= 488;
      opCodes[4084] <= 488;
      opCodes[4087] <= 488;
      opCodes[4148] <= 488;
      opCodes[4151] <= 488;
      opCodes[4189] <= 488;
      opCodes[4192] <= 488;
      opCodes[4230] <= 488;
      opCodes[4233] <= 488;
      opCodes[4271] <= 488;
      opCodes[4274] <= 488;
      opCodes[4312] <= 488;
      opCodes[4315] <= 488;
      opCodes[4353] <= 488;
      opCodes[4356] <= 488;
      opCodes[4394] <= 488;
      opCodes[4397] <= 488;
      opCodes[4435] <= 488;
      opCodes[4438] <= 488;
      opCodes[4476] <= 488;
      opCodes[4479] <= 488;
      opCodes[3715] <= 489;
      opCodes[3756] <= 489;
      opCodes[3797] <= 489;
      opCodes[3838] <= 489;
      opCodes[3879] <= 489;
      opCodes[3920] <= 489;
      opCodes[3961] <= 489;
      opCodes[4002] <= 489;
      opCodes[4085] <= 489;
      opCodes[4149] <= 489;
      opCodes[4190] <= 489;
      opCodes[4231] <= 489;
      opCodes[4272] <= 489;
      opCodes[4313] <= 489;
      opCodes[4354] <= 489;
      opCodes[4395] <= 489;
      opCodes[4436] <= 489;
      opCodes[4477] <= 489;
      opCodes[3718] <= 490;
      opCodes[3759] <= 490;
      opCodes[3800] <= 490;
      opCodes[3841] <= 490;
      opCodes[3882] <= 490;
      opCodes[3923] <= 490;
      opCodes[3964] <= 490;
      opCodes[4005] <= 490;
      opCodes[4088] <= 490;
      opCodes[4152] <= 490;
      opCodes[4193] <= 490;
      opCodes[4234] <= 490;
      opCodes[4275] <= 490;
      opCodes[4316] <= 490;
      opCodes[4357] <= 490;
      opCodes[4398] <= 490;
      opCodes[4439] <= 490;
      opCodes[4480] <= 490;
      opCodes[3719] <= 491;
      opCodes[3760] <= 491;
      opCodes[3801] <= 491;
      opCodes[3842] <= 491;
      opCodes[3883] <= 491;
      opCodes[3924] <= 491;
      opCodes[3965] <= 491;
      opCodes[4006] <= 491;
      opCodes[4089] <= 491;
      opCodes[4153] <= 491;
      opCodes[4194] <= 491;
      opCodes[4235] <= 491;
      opCodes[4276] <= 491;
      opCodes[4317] <= 491;
      opCodes[4358] <= 491;
      opCodes[4399] <= 491;
      opCodes[4440] <= 491;
      opCodes[4481] <= 491;
      opCodes[3720] <= 492;
      opCodes[3761] <= 492;
      opCodes[3802] <= 492;
      opCodes[3843] <= 492;
      opCodes[3884] <= 492;
      opCodes[3925] <= 492;
      opCodes[3966] <= 492;
      opCodes[4007] <= 492;
      opCodes[4090] <= 492;
      opCodes[4154] <= 492;
      opCodes[4195] <= 492;
      opCodes[4236] <= 492;
      opCodes[4277] <= 492;
      opCodes[4318] <= 492;
      opCodes[4359] <= 492;
      opCodes[4400] <= 492;
      opCodes[4441] <= 492;
      opCodes[4482] <= 492;
      opCodes[3721] <= 493;
      opCodes[3762] <= 493;
      opCodes[3803] <= 493;
      opCodes[3844] <= 493;
      opCodes[3885] <= 493;
      opCodes[3926] <= 493;
      opCodes[3967] <= 493;
      opCodes[4008] <= 493;
      opCodes[4091] <= 493;
      opCodes[4155] <= 493;
      opCodes[4196] <= 493;
      opCodes[4237] <= 493;
      opCodes[4278] <= 493;
      opCodes[4319] <= 493;
      opCodes[4360] <= 493;
      opCodes[4401] <= 493;
      opCodes[4442] <= 493;
      opCodes[4483] <= 493;
      opCodes[3725] <= 494;
      opCodes[3753] <= 495;
      opCodes[3766] <= 496;
      opCodes[3794] <= 497;
      opCodes[3807] <= 498;
      opCodes[3835] <= 499;
      opCodes[3848] <= 500;
      opCodes[3876] <= 501;
      opCodes[3889] <= 502;
      opCodes[3917] <= 503;
      opCodes[3930] <= 504;
      opCodes[3958] <= 505;
      opCodes[3971] <= 506;
      opCodes[3999] <= 507;
      opCodes[4012] <= 508;
      opCodes[4022] <= 509;
      opCodes[4050] <= 510;
      opCodes[4063] <= 511;
      opCodes[4077] <= 512;
      opCodes[4082] <= 513;
      opCodes[4095] <= 514;
      opCodes[4129] <= 515;
      opCodes[4170] <= 515;
      opCodes[4211] <= 515;
      opCodes[4252] <= 515;
      opCodes[4293] <= 515;
      opCodes[4334] <= 515;
      opCodes[4375] <= 515;
      opCodes[4416] <= 515;
      opCodes[4457] <= 515;
      opCodes[4146] <= 516;
      opCodes[4159] <= 517;
      opCodes[4187] <= 518;
      opCodes[4200] <= 519;
      opCodes[4228] <= 520;
      opCodes[4241] <= 521;
      opCodes[4269] <= 522;
      opCodes[4282] <= 523;
      opCodes[4310] <= 524;
      opCodes[4323] <= 525;
      opCodes[4351] <= 526;
      opCodes[4364] <= 527;
      opCodes[4392] <= 528;
      opCodes[4405] <= 529;
      opCodes[4433] <= 530;
      opCodes[4446] <= 531;
      opCodes[4474] <= 532;
      opCodes[4487] <= 533;
      opCodes[4497] <= 534;
      opCodes[4498] <= 535;
      opCodes[4499] <= 536;
      opCodes[4521] <= 537;
      opCodes[4532] <= 538;
      opCodes[5464] <= 538;
      opCodes[4534] <= 539;
      opCodes[4552] <= 539;
      opCodes[5466] <= 539;
      opCodes[5484] <= 539;
      opCodes[4535] <= 540;
      opCodes[4550] <= 540;
      opCodes[5467] <= 540;
      opCodes[5482] <= 540;
      opCodes[4536] <= 541;
      opCodes[4539] <= 541;
      opCodes[4555] <= 541;
      opCodes[5468] <= 541;
      opCodes[5471] <= 541;
      opCodes[5487] <= 541;
      opCodes[4537] <= 542;
      opCodes[4553] <= 542;
      opCodes[5469] <= 542;
      opCodes[5485] <= 542;
      opCodes[4544] <= 543;
      opCodes[5476] <= 543;
      opCodes[4545] <= 544;
      opCodes[4546] <= 545;
      opCodes[5478] <= 545;
      opCodes[4547] <= 546;
      opCodes[5479] <= 546;
      opCodes[4548] <= 547;
      opCodes[5480] <= 547;
      opCodes[4549] <= 548;
      opCodes[5481] <= 548;
      opCodes[4556] <= 549;
      opCodes[4560] <= 550;
      opCodes[4561] <= 551;
      opCodes[4562] <= 552;
      opCodes[4565] <= 553;
      opCodes[5495] <= 553;
      opCodes[4567] <= 554;
      opCodes[4569] <= 555;
      opCodes[4570] <= 556;
      opCodes[4571] <= 557;
      opCodes[4572] <= 558;
      opCodes[4575] <= 558;
      opCodes[4573] <= 559;
      opCodes[4576] <= 560;
      opCodes[4577] <= 561;
      opCodes[4578] <= 562;
      opCodes[4599] <= 562;
      opCodes[5001] <= 562;
      opCodes[5426] <= 562;
      opCodes[4580] <= 563;
      opCodes[4588] <= 563;
      opCodes[5003] <= 563;
      opCodes[5428] <= 563;
      opCodes[5439] <= 563;
      opCodes[5447] <= 563;
      opCodes[5458] <= 563;
      opCodes[4587] <= 564;
      opCodes[4598] <= 565;
      opCodes[4608] <= 566;
      opCodes[4609] <= 567;
      opCodes[4660] <= 567;
      opCodes[4701] <= 567;
      opCodes[4742] <= 567;
      opCodes[4783] <= 567;
      opCodes[4824] <= 567;
      opCodes[4865] <= 567;
      opCodes[4906] <= 567;
      opCodes[4947] <= 567;
      opCodes[4960] <= 567;
      opCodes[4988] <= 567;
      opCodes[5009] <= 567;
      opCodes[5059] <= 567;
      opCodes[5100] <= 567;
      opCodes[5141] <= 567;
      opCodes[5182] <= 567;
      opCodes[5223] <= 567;
      opCodes[5264] <= 567;
      opCodes[5305] <= 567;
      opCodes[5346] <= 567;
      opCodes[5387] <= 567;
      opCodes[4614] <= 568;
      opCodes[4968] <= 568;
      opCodes[4615] <= 569;
      opCodes[4633] <= 569;
      opCodes[4674] <= 569;
      opCodes[4715] <= 569;
      opCodes[4756] <= 569;
      opCodes[4797] <= 569;
      opCodes[4838] <= 569;
      opCodes[4879] <= 569;
      opCodes[4920] <= 569;
      opCodes[4969] <= 569;
      opCodes[5032] <= 569;
      opCodes[5073] <= 569;
      opCodes[5114] <= 569;
      opCodes[5155] <= 569;
      opCodes[5196] <= 569;
      opCodes[5237] <= 569;
      opCodes[5278] <= 569;
      opCodes[5319] <= 569;
      opCodes[5360] <= 569;
      opCodes[5398] <= 569;
      opCodes[5424] <= 569;
      opCodes[4620] <= 570;
      opCodes[4977] <= 570;
      opCodes[4621] <= 571;
      opCodes[4978] <= 571;
      opCodes[5013] <= 571;
      opCodes[4622] <= 572;
      opCodes[4624] <= 572;
      opCodes[4979] <= 572;
      opCodes[4982] <= 572;
      opCodes[4984] <= 572;
      opCodes[4623] <= 573;
      opCodes[4983] <= 573;
      opCodes[4625] <= 574;
      opCodes[4980] <= 574;
      opCodes[4985] <= 574;
      opCodes[4627] <= 575;
      opCodes[4987] <= 575;
      opCodes[4628] <= 576;
      opCodes[4629] <= 577;
      opCodes[5025] <= 577;
      opCodes[5028] <= 577;
      opCodes[4630] <= 578;
      opCodes[4671] <= 578;
      opCodes[4712] <= 578;
      opCodes[4753] <= 578;
      opCodes[4794] <= 578;
      opCodes[4835] <= 578;
      opCodes[4876] <= 578;
      opCodes[4917] <= 578;
      opCodes[5026] <= 578;
      opCodes[5029] <= 578;
      opCodes[5070] <= 578;
      opCodes[5111] <= 578;
      opCodes[5152] <= 578;
      opCodes[5193] <= 578;
      opCodes[5234] <= 578;
      opCodes[5275] <= 578;
      opCodes[5316] <= 578;
      opCodes[5357] <= 578;
      opCodes[4632] <= 579;
      opCodes[4673] <= 579;
      opCodes[4714] <= 579;
      opCodes[4755] <= 579;
      opCodes[4796] <= 579;
      opCodes[4837] <= 579;
      opCodes[4878] <= 579;
      opCodes[4919] <= 579;
      opCodes[4645] <= 580;
      opCodes[4656] <= 581;
      opCodes[4686] <= 582;
      opCodes[4697] <= 583;
      opCodes[4727] <= 584;
      opCodes[4738] <= 585;
      opCodes[4768] <= 586;
      opCodes[4779] <= 587;
      opCodes[4809] <= 588;
      opCodes[4820] <= 589;
      opCodes[4850] <= 590;
      opCodes[4861] <= 591;
      opCodes[4891] <= 592;
      opCodes[4902] <= 593;
      opCodes[4932] <= 594;
      opCodes[4943] <= 595;
      opCodes[4959] <= 596;
      opCodes[5000] <= 597;
      opCodes[5011] <= 598;
      opCodes[5020] <= 599;
      opCodes[5024] <= 600;
      opCodes[5031] <= 601;
      opCodes[5072] <= 601;
      opCodes[5113] <= 601;
      opCodes[5154] <= 601;
      opCodes[5195] <= 601;
      opCodes[5236] <= 601;
      opCodes[5277] <= 601;
      opCodes[5318] <= 601;
      opCodes[5359] <= 601;
      opCodes[5044] <= 602;
      opCodes[5055] <= 603;
      opCodes[5085] <= 604;
      opCodes[5096] <= 605;
      opCodes[5126] <= 606;
      opCodes[5137] <= 607;
      opCodes[5167] <= 608;
      opCodes[5178] <= 609;
      opCodes[5208] <= 610;
      opCodes[5219] <= 611;
      opCodes[5249] <= 612;
      opCodes[5260] <= 613;
      opCodes[5290] <= 614;
      opCodes[5301] <= 615;
      opCodes[5331] <= 616;
      opCodes[5342] <= 617;
      opCodes[5372] <= 618;
      opCodes[5383] <= 619;
      opCodes[5399] <= 620;
      opCodes[5400] <= 621;
      opCodes[5401] <= 622;
      opCodes[5423] <= 623;
      opCodes[5438] <= 624;
      opCodes[5445] <= 625;
      opCodes[5454] <= 626;
      opCodes[5477] <= 627;
      opCodes[5488] <= 628;
      opCodes[5492] <= 629;
      opCodes[5496] <= 630;
      opCodes[5499] <= 631;
      opCodes[5509] <= 632;
      opCodes[5522] <= 632;
      opCodes[5511] <= 633;
      opCodes[5517] <= 634;
      opCodes[5523] <= 635;
      opCodes[5530] <= 636;
      opCodes[5533] <= 636;
      opCodes[5532] <= 637;
      opCodes[5535] <= 638;
      opCodes[5536] <= 639;
      opCodes[5538] <= 640;
      opCodes[5553] <= 641;
      opCodes[5555] <= 642;
      opCodes[5557] <= 643;
      opCodes[5559] <= 644;
      opCodes[5561] <= 645;
      opCodes[5562] <= 646;
      opCodes[5590] <= 646;
      opCodes[5620] <= 646;
      opCodes[5658] <= 646;
      opCodes[5696] <= 646;
      opCodes[5734] <= 646;
      opCodes[5774] <= 646;
      opCodes[5791] <= 646;
      opCodes[5563] <= 647;
      opCodes[5565] <= 648;
      opCodes[5567] <= 649;
      opCodes[5568] <= 650;
      opCodes[5569] <= 651;
      opCodes[5593] <= 652;
      opCodes[5631] <= 652;
      opCodes[5669] <= 652;
      opCodes[5707] <= 652;
      opCodes[5745] <= 652;
      opCodes[5605] <= 653;
      opCodes[5616] <= 654;
      opCodes[5643] <= 655;
      opCodes[5654] <= 656;
      opCodes[5681] <= 657;
      opCodes[5692] <= 658;
      opCodes[5719] <= 659;
      opCodes[5730] <= 660;
      opCodes[5757] <= 661;
      opCodes[5768] <= 662;
      opCodes[5773] <= 663;
      opCodes[5787] <= 664;
      opCodes[5789] <= 665;
      opCodes[5793] <= 666;
      opCodes[5805] <= 667;
      opCodes[5816] <= 668;
      opCodes[5836] <= 669;
      opCodes[5849] <= 669;
      opCodes[5838] <= 670;
      opCodes[5844] <= 671;
      opCodes[5850] <= 672;
      opCodes[5858] <= 673;
      opCodes[5861] <= 674;
      opCodes[5864] <= 674;
      opCodes[5863] <= 675;
      opCodes[5866] <= 676;
      opCodes[5867] <= 677;

      $assignKey
      memory[183] <= 4; /* put data */
    end
    else begin                                                                  // Run
      //$display("%4d %4d %4d s=%4d f=%4d d=%4d", steps, step, intermediateValue, stop, found, data);
      case(opCodes[step])
           0 : begin intermediateValue <= memory[433]/*put_Key*/; /* get 1 */ step <= step + 1; end
           1 : begin memory[187]/*findAndInsert_Key*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
           2 : begin intermediateValue <= memory[432]/*put_Data*/; /* get 1 */ step <= step + 1; end
           3 : begin memory[186]/*findAndInsert_Data*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
           4 : begin intermediateValue <= memory[187]/*findAndInsert_Key*/; /* get 1 */ step <= step + 1; end
           5 : begin memory[189]/*find_Key*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
           6 : begin intermediateValue <= memory[217+memory[435]/*root*/]/*isLeaf[root]*/; /* get 2 */ step <= step + 1; end
           7 : begin memory[436]/*rootIsLeaf*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
           8 : begin intermediateValue <= memory[436]/*rootIsLeaf*/; /* get 1 */ step <= step + 1; end
           9 : begin if (intermediateValue == 0) step <=   44; else step = step + 1;/* endIfEq*/    end
          10 : begin memory[496]/*stuck*/ <= 0; /* set 1 */ step <= step + 1; end
          11 : begin intermediateValue <= memory[189]/*find_Key*/; /* get 1 */ step <= step + 1; end
          12 : begin memory[442]/*s_key*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          13 : begin memory[440]/*s_found*/ <= 0; /* set 1 */ step <= step + 1; end
          14 : begin memory[441]/*s_index*/ <= 0; /* set 1 */ step <= step + 1; end
          15 : begin intermediateValue <= memory[5+memory[496]/*stuck*/]/*current_size[stuck]*/; /* get 2 */ step <= step + 1; end
          16 : begin memory[492]/*stuckSearch_N*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          17 : begin intermediateValue <= memory[441]/*s_index*/ < memory[492]/*stuckSearch_N*/ ? -1 : memory[441]/*s_index*/ == memory[492]/*stuckSearch_N*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
          18 : begin if (intermediateValue >= 0) step <=   33; else step = step + 1;/* endIfGe*/    end
          19 : begin intermediateValue <= memory[442]/*s_key*/ < memory[234+memory[496]/*stuck*/*10+memory[441]/*s_index*/]/*keys[s_index,stuck]*/ ? -1 : memory[442]/*s_key*/ == memory[234+memory[496]/*stuck*/*10+memory[441]/*s_index*/]/*keys[s_index,stuck]*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
          20 : begin if (intermediateValue != 0) step <=   27; else step = step + 1;/* endIfNe*/    end
          21 : begin memory[440]/*s_found*/ <= 1; /* set 1 */ step <= step + 1; end
          22 : begin intermediateValue <= memory[234+memory[496]/*stuck*/*10+memory[441]/*s_index*/]/*keys[s_index,stuck]*/; /* get 3 */ step <= step + 1; end
          23 : begin intermediateValue <= memory[21+memory[496]/*stuck*/*10+memory[441]/*s_index*/]/*data[s_index,stuck]*/; /* get 3 */ step <= step + 1; end
          24 : begin memory[437]/*s_data*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          25 : begin step <=   33; /* end */ end
          26 : begin intermediateValue <= memory[441]/*s_index*/; /* get 1 */ step <= step + 1; end
          27 : begin intermediateValue <= 1 + intermediateValue;  /* add 1 */ step <= step + 1; end
          28 : begin memory[441]/*s_index*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          29 : begin step <= 17; /* start */ end
          30 : begin intermediateValue <= memory[435]/*root*/; /* get 1 */ step <= step + 1; end
          31 : begin memory[194]/*f_leaf*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          32 : begin intermediateValue <= memory[440]/*s_found*/; /* get 1 */ step <= step + 1; end
          33 : begin memory[184]/*f_found*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          34 : begin memory[188]/*f_index*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          35 : begin intermediateValue <= memory[442]/*s_key*/; /* get 1 */ step <= step + 1; end
          36 : begin memory[193]/*f_key*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          37 : begin intermediateValue <= memory[437]/*s_data*/; /* get 1 */ step <= step + 1; end
          38 : begin memory[183]/*f_data*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          39 : begin step <=   133; /* end */ end
          40 : begin memory[431]/*parent*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          41 : begin memory[190] <= 0; /* clear 1 */ step <= step + 1; end
          42 : begin intermediateValue <= memory[431]/*parent*/; /* get 1 */ step <= step + 1; end
          43 : begin memory[496]/*stuck*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          44 : begin intermediateValue <= memory[492]/*stuckSearch_N*/; /* get 1 */ step <= step + 1; end
          45 : begin intermediateValue <= -1 + intermediateValue;  /* add 1 */ step <= step + 1; end
          46 : begin if (intermediateValue >= 0) step <=   74; else step = step + 1;/* endIfGe*/    end
          47 : begin if (intermediateValue >  0) step <=   68; else step = step + 1;/* endIfGt*/    end
          48 : begin step <=   74; /* end */ end
          49 : begin step <= 58; /* start */ end
          50 : begin memory[4]/*child*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          51 : begin intermediateValue <= memory[4]/*child*/; /* get 1 */ step <= step + 1; end
          52 : begin memory[214]/*isALeaf*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          53 : begin intermediateValue <= memory[217+memory[214]/*isALeaf*/]/*isLeaf[isALeaf]*/; /* get 2 */ step <= step + 1; end
          54 : begin intermediateValue <= memory[214]/*isALeaf*/; /* get 1 */ step <= step + 1; end
          55 : begin if (intermediateValue == 0) step <=   123; else step = step + 1;/* endIfEq*/    end
          56 : begin if (intermediateValue >= 0) step <=   110; else step = step + 1;/* endIfGe*/    end
          57 : begin if (intermediateValue != 0) step <=   104; else step = step + 1;/* endIfNe*/    end
          58 : begin step <=   110; /* end */ end
          59 : begin step <= 94; /* start */ end
          60 : begin memory[191]/*find_result_leaf*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          61 : begin intermediateValue <= memory[191]/*find_result_leaf*/; /* get 1 */ step <= step + 1; end
          62 : begin intermediateValue <= memory[190]/*find_loop*/; /* get 1 */ step <= step + 1; end
          63 : begin memory[190]/*find_loop*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          64 : begin intermediateValue <= 9 <  intermediateValue ? -1 : 9 == intermediateValue ?  0 : +1; /* compare 1 */ step <= step + 1; end
          65 : begin if (intermediateValue >= 0) step <=   132; else step = step + 1;/* endIfGe*/    end
          66 : begin step <= 47; /* start */ end
          67 : begin stopped <= 1; end
          68 : begin intermediateValue <= memory[184]/*f_found*/; /* get 1 */ step <= step + 1; end
          69 : begin if (intermediateValue == 0) step <=   155; else step = step + 1;/* endIfEq*/    end
          70 : begin intermediateValue <= memory[194]/*f_leaf*/; /* get 1 */ step <= step + 1; end
          71 : begin intermediateValue <= memory[186]/*findAndInsert_Data*/; /* get 1 */ step <= step + 1; end
          72 : begin intermediateValue <= memory[188]/*f_index*/; /* get 1 */ step <= step + 1; end
          73 : begin memory[234+memory[496]/*stuck*/*10+memory[441]/*s_index*/]/*keys[s_index,stuck]*/ <= intermediateValue; /* set 3 */ step <= step + 1; end
          74 : begin memory[21+memory[496]/*stuck*/*10+memory[441]/*s_index*/]/*data[s_index,stuck]*/ <= intermediateValue; /* set 3 */ step <= step + 1; end
          75 : begin intermediateValue <= memory[441]/*s_index*/ < memory[5+memory[496]/*stuck*/]/*current_size[stuck]*/ ? -1 : memory[441]/*s_index*/ == memory[5+memory[496]/*stuck*/]/*current_size[stuck]*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
          76 : begin if (intermediateValue <  0) step <=   152; else step = step + 1;/* endIfLt*/    end
          77 : begin memory[5+memory[496]/*stuck*/]/*current_size[stuck]*/ <= intermediateValue; /* set 2 */ step <= step + 1; end
          78 : begin memory[212]/*f_success*/ <= 1; /* set 1 */ step <= step + 1; end
          79 : begin memory[192]/*f_inserted*/ <= 0; /* set 1 */ step <= step + 1; end
          80 : begin step <=   231; /* end */ end
          81 : begin memory[216]/*isFull*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          82 : begin intermediateValue <= memory[216]/*isFull*/; /* get 1 */ step <= step + 1; end
          83 : begin memory[394]/*leafSize*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          84 : begin intermediateValue <= memory[5+memory[394]/*leafSize*/]/*current_size[leafSize]*/; /* get 2 */ step <= step + 1; end
          85 : begin intermediateValue <= memory[394]/*leafSize*/; /* get 1 */ step <= step + 1; end
          86 : begin intermediateValue <= 8 <  intermediateValue ? -1 : 8 == intermediateValue ?  0 : +1; /* compare 1 */ step <= step + 1; end
          87 : begin intermediateValue <= intermediateValue >= 0 ? 1 : 0; /* ge */ step <= step + 1; end
          88 : begin if (intermediateValue >  0) step <=   229; else step = step + 1;/* endIfGt*/    end
          89 : begin if (intermediateValue >= 0) step <=   191; else step = step + 1;/* endIfGe*/    end
          90 : begin if (intermediateValue >  0) step <=   185; else step = step + 1;/* endIfGt*/    end
          91 : begin step <=   191; /* end */ end
          92 : begin step <= 175; /* start */ end
          93 : begin memory[488]/*stuckInsertElementAt_L*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          94 : begin memory[487]/*stuckInsertElementAt_i*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          95 : begin intermediateValue <= memory[487]/*stuckInsertElementAt_i*/; /* get 1 */ step <= step + 1; end
          96 : begin memory[486]/*stuckInsertElementAt_I*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
          97 : begin intermediateValue <= memory[486]/*stuckInsertElementAt_I*/; /* get 1 */ step <= step + 1; end
          98 : begin intermediateValue <= memory[487]/*stuckInsertElementAt_i*/ < memory[488]/*stuckInsertElementAt_L*/ ? -1 : memory[487]/*stuckInsertElementAt_i*/ == memory[488]/*stuckInsertElementAt_L*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
          99 : begin if (intermediateValue == 0) step <=   219; else step = step + 1;/* endIfEq*/    end
         100 : begin intermediateValue <= memory[234+memory[496]/*stuck*/*10+memory[486]/*stuckInsertElementAt_I*/]/*keys[stuckInsertElementAt_I,stuck]*/; /* get 3 */ step <= step + 1; end
         101 : begin memory[234+memory[496]/*stuck*/*10+memory[487]/*stuckInsertElementAt_i*/]/*keys[stuckInsertElementAt_i,stuck]*/ <= intermediateValue; /* set 3 */ step <= step + 1; end
         102 : begin intermediateValue <= memory[21+memory[496]/*stuck*/*10+memory[486]/*stuckInsertElementAt_I*/]/*data[stuckInsertElementAt_I,stuck]*/; /* get 3 */ step <= step + 1; end
         103 : begin memory[21+memory[496]/*stuck*/*10+memory[487]/*stuckInsertElementAt_i*/]/*data[stuckInsertElementAt_i,stuck]*/ <= intermediateValue; /* set 3 */ step <= step + 1; end
         104 : begin step <= 206; /* start */ end
         105 : begin memory[212]/*f_success*/ <= 0; /* set 1 */ step <= step + 1; end
         106 : begin intermediateValue <= memory[212]/*f_success*/; /* get 1 */ step <= step + 1; end
         107 : begin if (intermediateValue >  0) step <=   5869; else step = step + 1;/* endIfGt*/    end
         108 : begin memory[216] <= 0; /* clear 1 */ step <= step + 1; end
         109 : begin if (intermediateValue == 0) step <=   248; else step = step + 1;/* endIfEq*/    end
         110 : begin if (intermediateValue >  0) step <=   260; else step = step + 1;/* endIfGt*/    end
         111 : begin memory[3]/*branchSize*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         112 : begin intermediateValue <= memory[5+memory[3]/*branchSize*/]/*current_size[branchSize]*/; /* get 2 */ step <= step + 1; end
         113 : begin intermediateValue <= memory[3]/*branchSize*/; /* get 1 */ step <= step + 1; end
         114 : begin memory[215]/*isFullRoot*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         115 : begin intermediateValue <= memory[215]/*isFullRoot*/; /* get 1 */ step <= step + 1; end
         116 : begin if (intermediateValue == 0) step <=   1407; else step = step + 1;/* endIfEq*/    end
         117 : begin if (intermediateValue == 0) step <=   695; else step = step + 1;/* endIfEq*/    end
         118 : begin intermediateValue <= memory[195]/*freeChainHead*/; /* get 1 */ step <= step + 1; end
         119 : begin memory[462]/*splitLeafRoot_l*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         120 : begin intermediateValue <= memory[462]/*splitLeafRoot_l*/; /* get 1 */ step <= step + 1; end
         121 : begin if (intermediateValue >  0) step <=   273; else step = step + 1;/* endIfGt*/    end
         122 : begin intermediateValue <= memory[196+memory[462]/*splitLeafRoot_l*/]/*free[splitLeafRoot_l]*/; /* get 2 */ step <= step + 1; end
         123 : begin memory[195]/*freeChainHead*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         124 : begin memory[196+memory[462]/*splitLeafRoot_l*/]/*free[splitLeafRoot_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         125 : begin memory[217+memory[462]/*splitLeafRoot_l*/]/*isLeaf[splitLeafRoot_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         126 : begin memory[5+memory[462]/*splitLeafRoot_l*/]/*current_size[splitLeafRoot_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         127 : begin memory[234] <= 0; /* clear 2 */ step <= step + 1; end
         128 : begin memory[235] <= 0; /* clear 2 */ step <= step + 1; end
         129 : begin memory[236] <= 0; /* clear 2 */ step <= step + 1; end
         130 : begin memory[237] <= 0; /* clear 2 */ step <= step + 1; end
         131 : begin memory[238] <= 0; /* clear 2 */ step <= step + 1; end
         132 : begin memory[239] <= 0; /* clear 2 */ step <= step + 1; end
         133 : begin memory[240] <= 0; /* clear 2 */ step <= step + 1; end
         134 : begin memory[241] <= 0; /* clear 2 */ step <= step + 1; end
         135 : begin memory[242] <= 0; /* clear 2 */ step <= step + 1; end
         136 : begin memory[243] <= 0; /* clear 2 */ step <= step + 1; end
         137 : begin memory[21] <= 0; /* clear 2 */ step <= step + 1; end
         138 : begin memory[22] <= 0; /* clear 2 */ step <= step + 1; end
         139 : begin memory[23] <= 0; /* clear 2 */ step <= step + 1; end
         140 : begin memory[24] <= 0; /* clear 2 */ step <= step + 1; end
         141 : begin memory[25] <= 0; /* clear 2 */ step <= step + 1; end
         142 : begin memory[26] <= 0; /* clear 2 */ step <= step + 1; end
         143 : begin memory[27] <= 0; /* clear 2 */ step <= step + 1; end
         144 : begin memory[28] <= 0; /* clear 2 */ step <= step + 1; end
         145 : begin memory[29] <= 0; /* clear 2 */ step <= step + 1; end
         146 : begin memory[30] <= 0; /* clear 2 */ step <= step + 1; end
         147 : begin memory[439]/*setLeaf*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         148 : begin memory[217+memory[439]/*setLeaf*/]/*isLeaf[setLeaf]*/ <= 1; /* set 2 */ step <= step + 1; end
         149 : begin memory[463]/*splitLeafRoot_r*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         150 : begin intermediateValue <= memory[463]/*splitLeafRoot_r*/; /* get 1 */ step <= step + 1; end
         151 : begin if (intermediateValue >  0) step <=   306; else step = step + 1;/* endIfGt*/    end
         152 : begin intermediateValue <= memory[196+memory[463]/*splitLeafRoot_r*/]/*free[splitLeafRoot_r]*/; /* get 2 */ step <= step + 1; end
         153 : begin memory[196+memory[463]/*splitLeafRoot_r*/]/*free[splitLeafRoot_r]*/ <= 0; /* set 2 */ step <= step + 1; end
         154 : begin memory[217+memory[463]/*splitLeafRoot_r*/]/*isLeaf[splitLeafRoot_r]*/ <= 0; /* set 2 */ step <= step + 1; end
         155 : begin memory[5+memory[463]/*splitLeafRoot_r*/]/*current_size[splitLeafRoot_r]*/ <= 0; /* set 2 */ step <= step + 1; end
         156 : begin memory[441] <= 0; /* clear 1 */ step <= step + 1; end
         157 : begin memory[495]/*stuckShift_N*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         158 : begin memory[493]/*stuckShift_i*/ <= 0; /* set 1 */ step <= step + 1; end
         159 : begin memory[494]/*stuckShift_I*/ <= 1; /* set 1 */ step <= step + 1; end
         160 : begin intermediateValue <= memory[494]/*stuckShift_I*/ < memory[495]/*stuckShift_N*/ ? -1 : memory[494]/*stuckShift_I*/ == memory[495]/*stuckShift_N*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
         161 : begin if (intermediateValue >= 0) step <=   358; else step = step + 1;/* endIfGe*/    end
         162 : begin intermediateValue <= memory[234+memory[496]/*stuck*/*10+memory[494]/*stuckShift_I*/]/*keys[stuckShift_I,stuck]*/; /* get 3 */ step <= step + 1; end
         163 : begin memory[234+memory[496]/*stuck*/*10+memory[493]/*stuckShift_i*/]/*keys[stuckShift_i,stuck]*/ <= intermediateValue; /* set 3 */ step <= step + 1; end
         164 : begin intermediateValue <= memory[21+memory[496]/*stuck*/*10+memory[494]/*stuckShift_I*/]/*data[stuckShift_I,stuck]*/; /* get 3 */ step <= step + 1; end
         165 : begin memory[21+memory[496]/*stuck*/*10+memory[493]/*stuckShift_i*/]/*data[stuckShift_i,stuck]*/ <= intermediateValue; /* set 3 */ step <= step + 1; end
         166 : begin intermediateValue <= memory[493]/*stuckShift_i*/; /* get 1 */ step <= step + 1; end
         167 : begin memory[493]/*stuckShift_i*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         168 : begin intermediateValue <= memory[494]/*stuckShift_I*/; /* get 1 */ step <= step + 1; end
         169 : begin memory[494]/*stuckShift_I*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         170 : begin step <= 345; /* start */ end
         171 : begin if (intermediateValue >= 0) step <=   396; else step = step + 1;/* endIfGe*/    end
         172 : begin step <= 383; /* start */ end
         173 : begin if (intermediateValue >= 0) step <=   434; else step = step + 1;/* endIfGe*/    end
         174 : begin step <= 421; /* start */ end
         175 : begin if (intermediateValue >= 0) step <=   472; else step = step + 1;/* endIfGe*/    end
         176 : begin step <= 459; /* start */ end
         177 : begin if (intermediateValue >= 0) step <=   510; else step = step + 1;/* endIfGe*/    end
         178 : begin step <= 497; /* start */ end
         179 : begin if (intermediateValue >= 0) step <=   548; else step = step + 1;/* endIfGe*/    end
         180 : begin step <= 535; /* start */ end
         181 : begin if (intermediateValue >= 0) step <=   586; else step = step + 1;/* endIfGe*/    end
         182 : begin step <= 573; /* start */ end
         183 : begin if (intermediateValue >= 0) step <=   624; else step = step + 1;/* endIfGe*/    end
         184 : begin step <= 611; /* start */ end
         185 : begin memory[458]/*splitLeafRoot_first*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         186 : begin memory[461]/*splitLeafRoot_last*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         187 : begin intermediateValue <= memory[461]/*splitLeafRoot_last*/; /* get 1 */ step <= step + 1; end
         188 : begin memory[460]/*splitLeafRoot_kv*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         189 : begin intermediateValue <= memory[458]/*splitLeafRoot_first*/ + memory[460]/*splitLeafRoot_kv*/; /* add2 */ step <= step + 1; end
         190 : begin intermediateValue <= memory[460]/*splitLeafRoot_kv*/; /* get 1 */ step <= step + 1; end
         191 : begin intermediateValue <= intermediateValue >> 1; /* shift right */ step <= step + 1; end
         192 : begin memory[217+memory[435]/*root*/]/*isLeaf[root]*/ <= 0; /* set 2 */ step <= step + 1; end
         193 : begin memory[5+memory[496]/*stuck*/]/*current_size[stuck]*/ <= 0; /* set 2 */ step <= step + 1; end
         194 : begin if (intermediateValue >  0) step <=   1178; else step = step + 1;/* endIfGt*/    end
         195 : begin memory[448]/*splitBranchRoot_l*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         196 : begin intermediateValue <= memory[448]/*splitBranchRoot_l*/; /* get 1 */ step <= step + 1; end
         197 : begin if (intermediateValue >  0) step <=   702; else step = step + 1;/* endIfGt*/    end
         198 : begin intermediateValue <= memory[196+memory[448]/*splitBranchRoot_l*/]/*free[splitBranchRoot_l]*/; /* get 2 */ step <= step + 1; end
         199 : begin memory[196+memory[448]/*splitBranchRoot_l*/]/*free[splitBranchRoot_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         200 : begin memory[217+memory[448]/*splitBranchRoot_l*/]/*isLeaf[splitBranchRoot_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         201 : begin memory[5+memory[448]/*splitBranchRoot_l*/]/*current_size[splitBranchRoot_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         202 : begin memory[438]/*setBranch*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         203 : begin memory[217+memory[438]/*setBranch*/]/*isLeaf[setBranch]*/ <= 0; /* set 2 */ step <= step + 1; end
         204 : begin memory[450]/*splitBranchRoot_r*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         205 : begin intermediateValue <= memory[450]/*splitBranchRoot_r*/; /* get 1 */ step <= step + 1; end
         206 : begin if (intermediateValue >  0) step <=   735; else step = step + 1;/* endIfGt*/    end
         207 : begin intermediateValue <= memory[196+memory[450]/*splitBranchRoot_r*/]/*free[splitBranchRoot_r]*/; /* get 2 */ step <= step + 1; end
         208 : begin memory[196+memory[450]/*splitBranchRoot_r*/]/*free[splitBranchRoot_r]*/ <= 0; /* set 2 */ step <= step + 1; end
         209 : begin memory[217+memory[450]/*splitBranchRoot_r*/]/*isLeaf[splitBranchRoot_r]*/ <= 0; /* set 2 */ step <= step + 1; end
         210 : begin memory[5+memory[450]/*splitBranchRoot_r*/]/*current_size[splitBranchRoot_r]*/ <= 0; /* set 2 */ step <= step + 1; end
         211 : begin if (intermediateValue >= 0) step <=   787; else step = step + 1;/* endIfGe*/    end
         212 : begin step <= 774; /* start */ end
         213 : begin if (intermediateValue >= 0) step <=   825; else step = step + 1;/* endIfGe*/    end
         214 : begin step <= 812; /* start */ end
         215 : begin if (intermediateValue >= 0) step <=   863; else step = step + 1;/* endIfGe*/    end
         216 : begin step <= 850; /* start */ end
         217 : begin if (intermediateValue >= 0) step <=   901; else step = step + 1;/* endIfGe*/    end
         218 : begin step <= 888; /* start */ end
         219 : begin if (intermediateValue >= 0) step <=   939; else step = step + 1;/* endIfGe*/    end
         220 : begin step <= 926; /* start */ end
         221 : begin memory[449]/*splitBranchRoot_plk*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         222 : begin if (intermediateValue >= 0) step <=   981; else step = step + 1;/* endIfGe*/    end
         223 : begin step <= 968; /* start */ end
         224 : begin if (intermediateValue >= 0) step <=   1019; else step = step + 1;/* endIfGe*/    end
         225 : begin step <= 1006; /* start */ end
         226 : begin if (intermediateValue >= 0) step <=   1057; else step = step + 1;/* endIfGe*/    end
         227 : begin step <= 1044; /* start */ end
         228 : begin if (intermediateValue >= 0) step <=   1095; else step = step + 1;/* endIfGe*/    end
         229 : begin step <= 1082; /* start */ end
         230 : begin if (intermediateValue >= 0) step <=   1133; else step = step + 1;/* endIfGe*/    end
         231 : begin step <= 1120; /* start */ end
         232 : begin intermediateValue <= memory[449]/*splitBranchRoot_plk*/; /* get 1 */ step <= step + 1; end
         233 : begin if (intermediateValue == 0) step <=   1218; else step = step + 1;/* endIfEq*/    end
         234 : begin if (intermediateValue >= 0) step <=   1207; else step = step + 1;/* endIfGe*/    end
         235 : begin if (intermediateValue != 0) step <=   1201; else step = step + 1;/* endIfNe*/    end
         236 : begin step <=   1207; /* end */ end
         237 : begin step <= 1191; /* start */ end
         238 : begin step <=   1307; /* end */ end
         239 : begin if (intermediateValue >= 0) step <=   1248; else step = step + 1;/* endIfGe*/    end
         240 : begin if (intermediateValue >  0) step <=   1242; else step = step + 1;/* endIfGt*/    end
         241 : begin step <=   1248; /* end */ end
         242 : begin step <= 1232; /* start */ end
         243 : begin if (intermediateValue == 0) step <=   1297; else step = step + 1;/* endIfEq*/    end
         244 : begin if (intermediateValue >= 0) step <=   1284; else step = step + 1;/* endIfGe*/    end
         245 : begin if (intermediateValue != 0) step <=   1278; else step = step + 1;/* endIfNe*/    end
         246 : begin step <=   1284; /* end */ end
         247 : begin step <= 1268; /* start */ end
         248 : begin if (intermediateValue >= 0) step <=   1306; else step = step + 1;/* endIfGe*/    end
         249 : begin step <= 1221; /* start */ end
         250 : begin if (intermediateValue == 0) step <=   1329; else step = step + 1;/* endIfEq*/    end
         251 : begin if (intermediateValue <  0) step <=   1326; else step = step + 1;/* endIfLt*/    end
         252 : begin step <=   1405; /* end */ end
         253 : begin if (intermediateValue >  0) step <=   1403; else step = step + 1;/* endIfGt*/    end
         254 : begin if (intermediateValue >= 0) step <=   1365; else step = step + 1;/* endIfGe*/    end
         255 : begin if (intermediateValue >  0) step <=   1359; else step = step + 1;/* endIfGt*/    end
         256 : begin step <=   1365; /* end */ end
         257 : begin step <= 1349; /* start */ end
         258 : begin if (intermediateValue == 0) step <=   1393; else step = step + 1;/* endIfEq*/    end
         259 : begin step <= 1380; /* start */ end
         260 : begin memory[434] <= 0; /* clear 1 */ step <= step + 1; end
         261 : begin if (intermediateValue >= 0) step <=   1437; else step = step + 1;/* endIfGe*/    end
         262 : begin if (intermediateValue >  0) step <=   1431; else step = step + 1;/* endIfGt*/    end
         263 : begin step <=   1437; /* end */ end
         264 : begin step <= 1421; /* start */ end
         265 : begin if (intermediateValue == 0) step <=   5539; else step = step + 1;/* endIfEq*/    end
         266 : begin memory[456]/*splitLeaf_node*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         267 : begin memory[457]/*splitLeaf_parent*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         268 : begin memory[453]/*splitLeaf_index*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         269 : begin memory[455]/*splitLeaf_l*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         270 : begin intermediateValue <= memory[455]/*splitLeaf_l*/; /* get 1 */ step <= step + 1; end
         271 : begin if (intermediateValue >  0) step <=   1460; else step = step + 1;/* endIfGt*/    end
         272 : begin intermediateValue <= memory[196+memory[455]/*splitLeaf_l*/]/*free[splitLeaf_l]*/; /* get 2 */ step <= step + 1; end
         273 : begin memory[196+memory[455]/*splitLeaf_l*/]/*free[splitLeaf_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         274 : begin memory[217+memory[455]/*splitLeaf_l*/]/*isLeaf[splitLeaf_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         275 : begin memory[5+memory[455]/*splitLeaf_l*/]/*current_size[splitLeaf_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         276 : begin intermediateValue <= memory[456]/*splitLeaf_node*/; /* get 1 */ step <= step + 1; end
         277 : begin if (intermediateValue >= 0) step <=   1512; else step = step + 1;/* endIfGe*/    end
         278 : begin step <= 1499; /* start */ end
         279 : begin if (intermediateValue >= 0) step <=   1550; else step = step + 1;/* endIfGe*/    end
         280 : begin step <= 1537; /* start */ end
         281 : begin if (intermediateValue >= 0) step <=   1588; else step = step + 1;/* endIfGe*/    end
         282 : begin step <= 1575; /* start */ end
         283 : begin if (intermediateValue >= 0) step <=   1626; else step = step + 1;/* endIfGe*/    end
         284 : begin step <= 1613; /* start */ end
         285 : begin memory[451]/*splitLeaf_F*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         286 : begin memory[454]/*splitLeaf_L*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         287 : begin intermediateValue <= memory[451]/*splitLeaf_F*/; /* get 1 */ step <= step + 1; end
         288 : begin memory[452]/*splitLeaf_fl*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         289 : begin intermediateValue <= memory[454]/*splitLeaf_L*/ + memory[452]/*splitLeaf_fl*/; /* add2 */ step <= step + 1; end
         290 : begin intermediateValue <= memory[452]/*splitLeaf_fl*/; /* get 1 */ step <= step + 1; end
         291 : begin intermediateValue <= memory[457]/*splitLeaf_parent*/; /* get 1 */ step <= step + 1; end
         292 : begin intermediateValue <= memory[453]/*splitLeaf_index*/; /* get 1 */ step <= step + 1; end
         293 : begin if (intermediateValue == 0) step <=   1699; else step = step + 1;/* endIfEq*/    end
         294 : begin step <= 1686; /* start */ end
         295 : begin if (intermediateValue == 0) step <=   1746; else step = step + 1;/* endIfEq*/    end
         296 : begin if (intermediateValue >= 0) step <=   1735; else step = step + 1;/* endIfGe*/    end
         297 : begin if (intermediateValue != 0) step <=   1729; else step = step + 1;/* endIfNe*/    end
         298 : begin step <=   1735; /* end */ end
         299 : begin step <= 1719; /* start */ end
         300 : begin step <=   1835; /* end */ end
         301 : begin if (intermediateValue >= 0) step <=   1776; else step = step + 1;/* endIfGe*/    end
         302 : begin if (intermediateValue >  0) step <=   1770; else step = step + 1;/* endIfGt*/    end
         303 : begin step <=   1776; /* end */ end
         304 : begin step <= 1760; /* start */ end
         305 : begin if (intermediateValue == 0) step <=   1825; else step = step + 1;/* endIfEq*/    end
         306 : begin if (intermediateValue >= 0) step <=   1812; else step = step + 1;/* endIfGe*/    end
         307 : begin if (intermediateValue != 0) step <=   1806; else step = step + 1;/* endIfNe*/    end
         308 : begin step <=   1812; /* end */ end
         309 : begin step <= 1796; /* start */ end
         310 : begin if (intermediateValue >= 0) step <=   1834; else step = step + 1;/* endIfGe*/    end
         311 : begin step <= 1749; /* start */ end
         312 : begin if (intermediateValue == 0) step <=   1857; else step = step + 1;/* endIfEq*/    end
         313 : begin if (intermediateValue <  0) step <=   1854; else step = step + 1;/* endIfLt*/    end
         314 : begin step <=   1933; /* end */ end
         315 : begin if (intermediateValue >  0) step <=   1931; else step = step + 1;/* endIfGt*/    end
         316 : begin if (intermediateValue >= 0) step <=   1893; else step = step + 1;/* endIfGe*/    end
         317 : begin if (intermediateValue >  0) step <=   1887; else step = step + 1;/* endIfGt*/    end
         318 : begin step <=   1893; /* end */ end
         319 : begin step <= 1877; /* start */ end
         320 : begin if (intermediateValue == 0) step <=   1921; else step = step + 1;/* endIfEq*/    end
         321 : begin step <= 1908; /* start */ end
         322 : begin memory[397]/*merge_Key*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         323 : begin if (intermediateValue >  0) step <=   3598; else step = step + 1;/* endIfGt*/    end
         324 : begin memory[3] <= 0; /* clear 1 */ step <= step + 1; end
         325 : begin memory[427]/*mergeRoot_nP*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         326 : begin intermediateValue <= memory[427]/*mergeRoot_nP*/; /* get 1 */ step <= step + 1; end
         327 : begin intermediateValue <= 1 <  intermediateValue ? -1 : 1 == intermediateValue ?  0 : +1; /* compare 1 */ step <= step + 1; end
         328 : begin memory[424]/*mergeRoot_l*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         329 : begin memory[430]/*mergeRoot_r*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         330 : begin memory[213]/*hasLeavesForChildren*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         331 : begin intermediateValue <= memory[21+memory[213]/*hasLeavesForChildren*/*10+memory[0]]/*data[0,hasLeavesForChildren]*/; /* get 3 */ step <= step + 1; end
         332 : begin intermediateValue <= memory[213]/*hasLeavesForChildren*/; /* get 1 */ step <= step + 1; end
         333 : begin if (intermediateValue == 0) step <=   2716; else step = step + 1;/* endIfEq*/    end
         334 : begin intermediateValue <= memory[424]/*mergeRoot_l*/; /* get 1 */ step <= step + 1; end
         335 : begin memory[425]/*mergeRoot_nl*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         336 : begin intermediateValue <= memory[430]/*mergeRoot_r*/; /* get 1 */ step <= step + 1; end
         337 : begin memory[428]/*mergeRoot_nr*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         338 : begin intermediateValue <= memory[425]/*mergeRoot_nl*/; /* get 1 */ step <= step + 1; end
         339 : begin memory[426]/*mergeRoot_nlr*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         340 : begin intermediateValue <= memory[428]/*mergeRoot_nr*/ + memory[426]/*mergeRoot_nlr*/; /* add2 */ step <= step + 1; end
         341 : begin intermediateValue <= memory[426]/*mergeRoot_nlr*/; /* get 1 */ step <= step + 1; end
         342 : begin intermediateValue <= 0 <  intermediateValue ? -1 : 0 == intermediateValue ?  0 : +1; /* compare 1 */ step <= step + 1; end
         343 : begin if (intermediateValue <= 0) step <=   2329; else step = step + 1;/* endIfLe*/    end
         344 : begin if (intermediateValue >= 0) step <=   2028; else step = step + 1;/* endIfGe*/    end
         345 : begin step <= 2015; /* start */ end
         346 : begin if (intermediateValue >= 0) step <=   2069; else step = step + 1;/* endIfGe*/    end
         347 : begin step <= 2056; /* start */ end
         348 : begin intermediateValue <= 2 <  intermediateValue ? -1 : 2 == intermediateValue ?  0 : +1; /* compare 1 */ step <= step + 1; end
         349 : begin if (intermediateValue >= 0) step <=   2110; else step = step + 1;/* endIfGe*/    end
         350 : begin step <= 2097; /* start */ end
         351 : begin intermediateValue <= 3 <  intermediateValue ? -1 : 3 == intermediateValue ?  0 : +1; /* compare 1 */ step <= step + 1; end
         352 : begin if (intermediateValue >= 0) step <=   2151; else step = step + 1;/* endIfGe*/    end
         353 : begin step <= 2138; /* start */ end
         354 : begin intermediateValue <= 4 <  intermediateValue ? -1 : 4 == intermediateValue ?  0 : +1; /* compare 1 */ step <= step + 1; end
         355 : begin if (intermediateValue >= 0) step <=   2192; else step = step + 1;/* endIfGe*/    end
         356 : begin step <= 2179; /* start */ end
         357 : begin intermediateValue <= 5 <  intermediateValue ? -1 : 5 == intermediateValue ?  0 : +1; /* compare 1 */ step <= step + 1; end
         358 : begin if (intermediateValue >= 0) step <=   2233; else step = step + 1;/* endIfGe*/    end
         359 : begin step <= 2220; /* start */ end
         360 : begin intermediateValue <= 6 <  intermediateValue ? -1 : 6 == intermediateValue ?  0 : +1; /* compare 1 */ step <= step + 1; end
         361 : begin if (intermediateValue >= 0) step <=   2274; else step = step + 1;/* endIfGe*/    end
         362 : begin step <= 2261; /* start */ end
         363 : begin intermediateValue <= 7 <  intermediateValue ? -1 : 7 == intermediateValue ?  0 : +1; /* compare 1 */ step <= step + 1; end
         364 : begin if (intermediateValue >= 0) step <=   2315; else step = step + 1;/* endIfGe*/    end
         365 : begin step <= 2302; /* start */ end
         366 : begin intermediateValue <= memory[428]/*mergeRoot_nr*/; /* get 1 */ step <= step + 1; end
         367 : begin if (intermediateValue <= 0) step <=   2657; else step = step + 1;/* endIfLe*/    end
         368 : begin if (intermediateValue >= 0) step <=   2356; else step = step + 1;/* endIfGe*/    end
         369 : begin step <= 2343; /* start */ end
         370 : begin if (intermediateValue >= 0) step <=   2397; else step = step + 1;/* endIfGe*/    end
         371 : begin step <= 2384; /* start */ end
         372 : begin if (intermediateValue >= 0) step <=   2438; else step = step + 1;/* endIfGe*/    end
         373 : begin step <= 2425; /* start */ end
         374 : begin if (intermediateValue >= 0) step <=   2479; else step = step + 1;/* endIfGe*/    end
         375 : begin step <= 2466; /* start */ end
         376 : begin if (intermediateValue >= 0) step <=   2520; else step = step + 1;/* endIfGe*/    end
         377 : begin step <= 2507; /* start */ end
         378 : begin if (intermediateValue >= 0) step <=   2561; else step = step + 1;/* endIfGe*/    end
         379 : begin step <= 2548; /* start */ end
         380 : begin if (intermediateValue >= 0) step <=   2602; else step = step + 1;/* endIfGe*/    end
         381 : begin step <= 2589; /* start */ end
         382 : begin if (intermediateValue >= 0) step <=   2643; else step = step + 1;/* endIfGe*/    end
         383 : begin step <= 2630; /* start */ end
         384 : begin memory[196+memory[424]/*mergeRoot_l*/]/*free[mergeRoot_l]*/ <= -1; /* set 2 */ step <= step + 1; end
         385 : begin memory[217+memory[424]/*mergeRoot_l*/]/*isLeaf[mergeRoot_l]*/ <= -1; /* set 2 */ step <= step + 1; end
         386 : begin memory[5+memory[424]/*mergeRoot_l*/]/*current_size[mergeRoot_l]*/ <= -1; /* set 2 */ step <= step + 1; end
         387 : begin memory[234] <= -1; /* clear 2 */ step <= step + 1; end
         388 : begin memory[235] <= -1; /* clear 2 */ step <= step + 1; end
         389 : begin memory[236] <= -1; /* clear 2 */ step <= step + 1; end
         390 : begin memory[237] <= -1; /* clear 2 */ step <= step + 1; end
         391 : begin memory[238] <= -1; /* clear 2 */ step <= step + 1; end
         392 : begin memory[239] <= -1; /* clear 2 */ step <= step + 1; end
         393 : begin memory[240] <= -1; /* clear 2 */ step <= step + 1; end
         394 : begin memory[241] <= -1; /* clear 2 */ step <= step + 1; end
         395 : begin memory[242] <= -1; /* clear 2 */ step <= step + 1; end
         396 : begin memory[243] <= -1; /* clear 2 */ step <= step + 1; end
         397 : begin memory[21] <= -1; /* clear 2 */ step <= step + 1; end
         398 : begin memory[22] <= -1; /* clear 2 */ step <= step + 1; end
         399 : begin memory[23] <= -1; /* clear 2 */ step <= step + 1; end
         400 : begin memory[24] <= -1; /* clear 2 */ step <= step + 1; end
         401 : begin memory[25] <= -1; /* clear 2 */ step <= step + 1; end
         402 : begin memory[26] <= -1; /* clear 2 */ step <= step + 1; end
         403 : begin memory[27] <= -1; /* clear 2 */ step <= step + 1; end
         404 : begin memory[28] <= -1; /* clear 2 */ step <= step + 1; end
         405 : begin memory[29] <= -1; /* clear 2 */ step <= step + 1; end
         406 : begin memory[30] <= -1; /* clear 2 */ step <= step + 1; end
         407 : begin memory[196+memory[424]/*mergeRoot_l*/]/*free[mergeRoot_l]*/ <= intermediateValue; /* set 2 */ step <= step + 1; end
         408 : begin memory[196+memory[430]/*mergeRoot_r*/]/*free[mergeRoot_r]*/ <= -1; /* set 2 */ step <= step + 1; end
         409 : begin memory[217+memory[430]/*mergeRoot_r*/]/*isLeaf[mergeRoot_r]*/ <= -1; /* set 2 */ step <= step + 1; end
         410 : begin memory[5+memory[430]/*mergeRoot_r*/]/*current_size[mergeRoot_r]*/ <= -1; /* set 2 */ step <= step + 1; end
         411 : begin memory[196+memory[430]/*mergeRoot_r*/]/*free[mergeRoot_r]*/ <= intermediateValue; /* set 2 */ step <= step + 1; end
         412 : begin memory[429]/*mergeRoot_pkn*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         413 : begin if (intermediateValue <= 0) step <=   3125; else step = step + 1;/* endIfLe*/    end
         414 : begin if (intermediateValue >= 0) step <=   2783; else step = step + 1;/* endIfGe*/    end
         415 : begin step <= 2770; /* start */ end
         416 : begin if (intermediateValue >= 0) step <=   2824; else step = step + 1;/* endIfGe*/    end
         417 : begin step <= 2811; /* start */ end
         418 : begin if (intermediateValue >= 0) step <=   2865; else step = step + 1;/* endIfGe*/    end
         419 : begin step <= 2852; /* start */ end
         420 : begin if (intermediateValue >= 0) step <=   2906; else step = step + 1;/* endIfGe*/    end
         421 : begin step <= 2893; /* start */ end
         422 : begin if (intermediateValue >= 0) step <=   2947; else step = step + 1;/* endIfGe*/    end
         423 : begin step <= 2934; /* start */ end
         424 : begin if (intermediateValue >= 0) step <=   2988; else step = step + 1;/* endIfGe*/    end
         425 : begin step <= 2975; /* start */ end
         426 : begin if (intermediateValue >= 0) step <=   3029; else step = step + 1;/* endIfGe*/    end
         427 : begin step <= 3016; /* start */ end
         428 : begin if (intermediateValue >= 0) step <=   3070; else step = step + 1;/* endIfGe*/    end
         429 : begin step <= 3057; /* start */ end
         430 : begin if (intermediateValue >= 0) step <=   3111; else step = step + 1;/* endIfGe*/    end
         431 : begin step <= 3098; /* start */ end
         432 : begin intermediateValue <= memory[429]/*mergeRoot_pkn*/; /* get 1 */ step <= step + 1; end
         433 : begin if (intermediateValue <= 0) step <=   3518; else step = step + 1;/* endIfLe*/    end
         434 : begin if (intermediateValue >= 0) step <=   3176; else step = step + 1;/* endIfGe*/    end
         435 : begin step <= 3163; /* start */ end
         436 : begin if (intermediateValue >= 0) step <=   3217; else step = step + 1;/* endIfGe*/    end
         437 : begin step <= 3204; /* start */ end
         438 : begin if (intermediateValue >= 0) step <=   3258; else step = step + 1;/* endIfGe*/    end
         439 : begin step <= 3245; /* start */ end
         440 : begin if (intermediateValue >= 0) step <=   3299; else step = step + 1;/* endIfGe*/    end
         441 : begin step <= 3286; /* start */ end
         442 : begin if (intermediateValue >= 0) step <=   3340; else step = step + 1;/* endIfGe*/    end
         443 : begin step <= 3327; /* start */ end
         444 : begin if (intermediateValue >= 0) step <=   3381; else step = step + 1;/* endIfGe*/    end
         445 : begin step <= 3368; /* start */ end
         446 : begin if (intermediateValue >= 0) step <=   3422; else step = step + 1;/* endIfGe*/    end
         447 : begin step <= 3409; /* start */ end
         448 : begin if (intermediateValue >= 0) step <=   3463; else step = step + 1;/* endIfGe*/    end
         449 : begin step <= 3450; /* start */ end
         450 : begin if (intermediateValue >= 0) step <=   3504; else step = step + 1;/* endIfGe*/    end
         451 : begin step <= 3491; /* start */ end
         452 : begin memory[409] <= 0; /* clear 1 */ step <= step + 1; end
         453 : begin memory[409]/*merge_loop*/ <= 0; /* set 1 */ step <= step + 1; end
         454 : begin if (intermediateValue >  0) step <=   5538; else step = step + 1;/* endIfGt*/    end
         455 : begin memory[395]/*merge_indexLimit*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         456 : begin intermediateValue <= memory[395]/*merge_indexLimit*/; /* get 1 */ step <= step + 1; end
         457 : begin memory[396]/*merge_indices*/ <= 0; /* set 1 */ step <= step + 1; end
         458 : begin intermediateValue <= memory[396]/*merge_indices*/ < memory[395]/*merge_indexLimit*/ ? -1 : memory[396]/*merge_indices*/ == memory[395]/*merge_indexLimit*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
         459 : begin if (intermediateValue >= 0) step <=   5497; else step = step + 1;/* endIfGe*/    end
         460 : begin memory[404]/*mergeLeftSibling_parent*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         461 : begin intermediateValue <= memory[396]/*merge_indices*/; /* get 1 */ step <= step + 1; end
         462 : begin memory[399]/*mergeLeftSibling_index*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         463 : begin memory[408] <= 0; /* clear 1 */ step <= step + 1; end
         464 : begin intermediateValue <= memory[399]/*mergeLeftSibling_index*/; /* get 1 */ step <= step + 1; end
         465 : begin if (intermediateValue == 0) step <=   4561; else step = step + 1;/* endIfEq*/    end
         466 : begin intermediateValue <= memory[404]/*mergeLeftSibling_parent*/; /* get 1 */ step <= step + 1; end
         467 : begin memory[398]/*mergeLeftSibling_bs*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         468 : begin intermediateValue <= memory[399]/*mergeLeftSibling_index*/ < memory[398]/*mergeLeftSibling_bs*/ ? -1 : memory[399]/*mergeLeftSibling_index*/ == memory[398]/*mergeLeftSibling_bs*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
         469 : begin if (intermediateValue >= 0) step <=   4561; else step = step + 1;/* endIfGe*/    end
         470 : begin memory[400]/*mergeLeftSibling_l*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         471 : begin memory[405]/*mergeLeftSibling_r*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         472 : begin if (intermediateValue == 0) step <=   4021; else step = step + 1;/* endIfEq*/    end
         473 : begin intermediateValue <= memory[400]/*mergeLeftSibling_l*/; /* get 1 */ step <= step + 1; end
         474 : begin memory[401]/*mergeLeftSibling_nl*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         475 : begin intermediateValue <= memory[405]/*mergeLeftSibling_r*/; /* get 1 */ step <= step + 1; end
         476 : begin memory[403]/*mergeLeftSibling_nr*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         477 : begin intermediateValue <= memory[401]/*mergeLeftSibling_nl*/; /* get 1 */ step <= step + 1; end
         478 : begin memory[402]/*mergeLeftSibling_nlr*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         479 : begin intermediateValue <= memory[403]/*mergeLeftSibling_nr*/ + memory[402]/*mergeLeftSibling_nlr*/; /* add2 */ step <= step + 1; end
         480 : begin intermediateValue <= memory[402]/*mergeLeftSibling_nlr*/; /* get 1 */ step <= step + 1; end
         481 : begin intermediateValue <= memory[5+memory[400]/*mergeLeftSibling_l*/]/*current_size[mergeLeftSibling_l]*/; /* get 2 */ step <= step + 1; end
         482 : begin memory[406]/*mergeLeftSibling_size*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         483 : begin intermediateValue <= memory[406]/*mergeLeftSibling_size*/; /* get 1 */ step <= step + 1; end
         484 : begin if (intermediateValue <= 0) step <=   4021; else step = step + 1;/* endIfLe*/    end
         485 : begin memory[497]/*stuckUnshift_i*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         486 : begin intermediateValue <= memory[497]/*stuckUnshift_i*/; /* get 1 */ step <= step + 1; end
         487 : begin if (intermediateValue <= 0) step <=   3726; else step = step + 1;/* endIfLe*/    end
         488 : begin memory[498]/*stuckUnshift_I*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         489 : begin intermediateValue <= memory[498]/*stuckUnshift_I*/; /* get 1 */ step <= step + 1; end
         490 : begin intermediateValue <= memory[234+memory[496]/*stuck*/*10+memory[498]/*stuckUnshift_I*/]/*keys[stuckUnshift_I,stuck]*/; /* get 3 */ step <= step + 1; end
         491 : begin memory[234+memory[496]/*stuck*/*10+memory[497]/*stuckUnshift_i*/]/*keys[stuckUnshift_i,stuck]*/ <= intermediateValue; /* set 3 */ step <= step + 1; end
         492 : begin intermediateValue <= memory[21+memory[496]/*stuck*/*10+memory[498]/*stuckUnshift_I*/]/*data[stuckUnshift_I,stuck]*/; /* get 3 */ step <= step + 1; end
         493 : begin memory[21+memory[496]/*stuck*/*10+memory[497]/*stuckUnshift_i*/]/*data[stuckUnshift_i,stuck]*/ <= intermediateValue; /* set 3 */ step <= step + 1; end
         494 : begin step <= 3711; /* start */ end
         495 : begin if (intermediateValue <= 0) step <=   3767; else step = step + 1;/* endIfLe*/    end
         496 : begin step <= 3752; /* start */ end
         497 : begin if (intermediateValue <= 0) step <=   3808; else step = step + 1;/* endIfLe*/    end
         498 : begin step <= 3793; /* start */ end
         499 : begin if (intermediateValue <= 0) step <=   3849; else step = step + 1;/* endIfLe*/    end
         500 : begin step <= 3834; /* start */ end
         501 : begin if (intermediateValue <= 0) step <=   3890; else step = step + 1;/* endIfLe*/    end
         502 : begin step <= 3875; /* start */ end
         503 : begin if (intermediateValue <= 0) step <=   3931; else step = step + 1;/* endIfLe*/    end
         504 : begin step <= 3916; /* start */ end
         505 : begin if (intermediateValue <= 0) step <=   3972; else step = step + 1;/* endIfLe*/    end
         506 : begin step <= 3957; /* start */ end
         507 : begin if (intermediateValue <= 0) step <=   4013; else step = step + 1;/* endIfLe*/    end
         508 : begin step <= 3998; /* start */ end
         509 : begin if (intermediateValue >  0) step <=   4496; else step = step + 1;/* endIfGt*/    end
         510 : begin if (intermediateValue >  0) step <=   4561; else step = step + 1;/* endIfGt*/    end
         511 : begin memory[407]/*mergeLeftSibling_t*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         512 : begin intermediateValue <= memory[407]/*mergeLeftSibling_t*/; /* get 1 */ step <= step + 1; end
         513 : begin if (intermediateValue <= 0) step <=   4096; else step = step + 1;/* endIfLe*/    end
         514 : begin step <= 4081; /* start */ end
         515 : begin if (intermediateValue <= 0) step <=   4496; else step = step + 1;/* endIfLe*/    end
         516 : begin if (intermediateValue <= 0) step <=   4160; else step = step + 1;/* endIfLe*/    end
         517 : begin step <= 4145; /* start */ end
         518 : begin if (intermediateValue <= 0) step <=   4201; else step = step + 1;/* endIfLe*/    end
         519 : begin step <= 4186; /* start */ end
         520 : begin if (intermediateValue <= 0) step <=   4242; else step = step + 1;/* endIfLe*/    end
         521 : begin step <= 4227; /* start */ end
         522 : begin if (intermediateValue <= 0) step <=   4283; else step = step + 1;/* endIfLe*/    end
         523 : begin step <= 4268; /* start */ end
         524 : begin if (intermediateValue <= 0) step <=   4324; else step = step + 1;/* endIfLe*/    end
         525 : begin step <= 4309; /* start */ end
         526 : begin if (intermediateValue <= 0) step <=   4365; else step = step + 1;/* endIfLe*/    end
         527 : begin step <= 4350; /* start */ end
         528 : begin if (intermediateValue <= 0) step <=   4406; else step = step + 1;/* endIfLe*/    end
         529 : begin step <= 4391; /* start */ end
         530 : begin if (intermediateValue <= 0) step <=   4447; else step = step + 1;/* endIfLe*/    end
         531 : begin step <= 4432; /* start */ end
         532 : begin if (intermediateValue <= 0) step <=   4488; else step = step + 1;/* endIfLe*/    end
         533 : begin step <= 4473; /* start */ end
         534 : begin memory[196+memory[400]/*mergeLeftSibling_l*/]/*free[mergeLeftSibling_l]*/ <= -1; /* set 2 */ step <= step + 1; end
         535 : begin memory[217+memory[400]/*mergeLeftSibling_l*/]/*isLeaf[mergeLeftSibling_l]*/ <= -1; /* set 2 */ step <= step + 1; end
         536 : begin memory[5+memory[400]/*mergeLeftSibling_l*/]/*current_size[mergeLeftSibling_l]*/ <= -1; /* set 2 */ step <= step + 1; end
         537 : begin memory[196+memory[400]/*mergeLeftSibling_l*/]/*free[mergeLeftSibling_l]*/ <= intermediateValue; /* set 2 */ step <= step + 1; end
         538 : begin memory[491]/*stuckRemoveElementAt_N*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         539 : begin memory[490]/*stuckRemoveElementAt_i*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         540 : begin intermediateValue <= memory[490]/*stuckRemoveElementAt_i*/; /* get 1 */ step <= step + 1; end
         541 : begin memory[489]/*stuckRemoveElementAt_I*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         542 : begin intermediateValue <= memory[489]/*stuckRemoveElementAt_I*/; /* get 1 */ step <= step + 1; end
         543 : begin intermediateValue <= memory[489]/*stuckRemoveElementAt_I*/ < memory[491]/*stuckRemoveElementAt_N*/ ? -1 : memory[489]/*stuckRemoveElementAt_I*/ == memory[491]/*stuckRemoveElementAt_N*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
         544 : begin if (intermediateValue == 0) step <=   4557; else step = step + 1;/* endIfEq*/    end
         545 : begin intermediateValue <= memory[234+memory[496]/*stuck*/*10+memory[489]/*stuckRemoveElementAt_I*/]/*keys[stuckRemoveElementAt_I,stuck]*/; /* get 3 */ step <= step + 1; end
         546 : begin memory[234+memory[496]/*stuck*/*10+memory[490]/*stuckRemoveElementAt_i*/]/*keys[stuckRemoveElementAt_i,stuck]*/ <= intermediateValue; /* set 3 */ step <= step + 1; end
         547 : begin intermediateValue <= memory[21+memory[496]/*stuck*/*10+memory[489]/*stuckRemoveElementAt_I*/]/*data[stuckRemoveElementAt_I,stuck]*/; /* get 3 */ step <= step + 1; end
         548 : begin memory[21+memory[496]/*stuck*/*10+memory[490]/*stuckRemoveElementAt_i*/]/*data[stuckRemoveElementAt_i,stuck]*/ <= intermediateValue; /* set 3 */ step <= step + 1; end
         549 : begin step <= 4544; /* start */ end
         550 : begin memory[408] <= 1; /* clear 1 */ step <= step + 1; end
         551 : begin intermediateValue <= memory[408]/*mergeLeftSibling*/; /* get 1 */ step <= step + 1; end
         552 : begin if (intermediateValue == 0) step <=   4566; else step = step + 1;/* endIfEq*/    end
         553 : begin memory[396]/*merge_indices*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         554 : begin memory[418]/*mergeRightSibling_parent*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         555 : begin memory[412]/*mergeRightSibling_index*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         556 : begin memory[423] <= 0; /* clear 1 */ step <= step + 1; end
         557 : begin intermediateValue <= memory[5+memory[418]/*mergeRightSibling_parent*/]/*current_size[mergeRightSibling_parent]*/; /* get 2 */ step <= step + 1; end
         558 : begin memory[410]/*mergeRightSibling_bs*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         559 : begin intermediateValue <= memory[410]/*mergeRightSibling_bs*/; /* get 1 */ step <= step + 1; end
         560 : begin intermediateValue <= memory[412]/*mergeRightSibling_index*/ < memory[410]/*mergeRightSibling_bs*/ ? -1 : memory[412]/*mergeRightSibling_index*/ == memory[410]/*mergeRightSibling_bs*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
         561 : begin if (intermediateValue >= 0) step <=   5493; else step = step + 1;/* endIfGe*/    end
         562 : begin intermediateValue <= memory[418]/*mergeRightSibling_parent*/; /* get 1 */ step <= step + 1; end
         563 : begin intermediateValue <= memory[412]/*mergeRightSibling_index*/; /* get 1 */ step <= step + 1; end
         564 : begin memory[414]/*mergeRightSibling_l*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         565 : begin memory[420]/*mergeRightSibling_r*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         566 : begin if (intermediateValue == 0) step <=   4958; else step = step + 1;/* endIfEq*/    end
         567 : begin intermediateValue <= memory[414]/*mergeRightSibling_l*/; /* get 1 */ step <= step + 1; end
         568 : begin memory[415]/*mergeRightSibling_nl*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         569 : begin intermediateValue <= memory[420]/*mergeRightSibling_r*/; /* get 1 */ step <= step + 1; end
         570 : begin memory[417]/*mergeRightSibling_nr*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         571 : begin intermediateValue <= memory[415]/*mergeRightSibling_nl*/; /* get 1 */ step <= step + 1; end
         572 : begin memory[416]/*mergeRightSibling_nlr*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         573 : begin intermediateValue <= memory[417]/*mergeRightSibling_nr*/ + memory[416]/*mergeRightSibling_nlr*/; /* add2 */ step <= step + 1; end
         574 : begin intermediateValue <= memory[416]/*mergeRightSibling_nlr*/; /* get 1 */ step <= step + 1; end
         575 : begin if (intermediateValue >  0) step <=   5493; else step = step + 1;/* endIfGt*/    end
         576 : begin intermediateValue <= memory[5+memory[420]/*mergeRightSibling_r*/]/*current_size[mergeRightSibling_r]*/; /* get 2 */ step <= step + 1; end
         577 : begin memory[421]/*mergeRightSibling_size*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         578 : begin intermediateValue <= memory[421]/*mergeRightSibling_size*/; /* get 1 */ step <= step + 1; end
         579 : begin if (intermediateValue <= 0) step <=   4958; else step = step + 1;/* endIfLe*/    end
         580 : begin if (intermediateValue >= 0) step <=   4657; else step = step + 1;/* endIfGe*/    end
         581 : begin step <= 4644; /* start */ end
         582 : begin if (intermediateValue >= 0) step <=   4698; else step = step + 1;/* endIfGe*/    end
         583 : begin step <= 4685; /* start */ end
         584 : begin if (intermediateValue >= 0) step <=   4739; else step = step + 1;/* endIfGe*/    end
         585 : begin step <= 4726; /* start */ end
         586 : begin if (intermediateValue >= 0) step <=   4780; else step = step + 1;/* endIfGe*/    end
         587 : begin step <= 4767; /* start */ end
         588 : begin if (intermediateValue >= 0) step <=   4821; else step = step + 1;/* endIfGe*/    end
         589 : begin step <= 4808; /* start */ end
         590 : begin if (intermediateValue >= 0) step <=   4862; else step = step + 1;/* endIfGe*/    end
         591 : begin step <= 4849; /* start */ end
         592 : begin if (intermediateValue >= 0) step <=   4903; else step = step + 1;/* endIfGe*/    end
         593 : begin step <= 4890; /* start */ end
         594 : begin if (intermediateValue >= 0) step <=   4944; else step = step + 1;/* endIfGe*/    end
         595 : begin step <= 4931; /* start */ end
         596 : begin if (intermediateValue >  0) step <=   5398; else step = step + 1;/* endIfGt*/    end
         597 : begin memory[413]/*mergeRightSibling_ld*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         598 : begin intermediateValue <= memory[413]/*mergeRightSibling_ld*/; /* get 1 */ step <= step + 1; end
         599 : begin if (intermediateValue <  0) step <=   5024; else step = step + 1;/* endIfLt*/    end
         600 : begin intermediateValue <= memory[417]/*mergeRightSibling_nr*/; /* get 1 */ step <= step + 1; end
         601 : begin if (intermediateValue <= 0) step <=   5398; else step = step + 1;/* endIfLe*/    end
         602 : begin if (intermediateValue >= 0) step <=   5056; else step = step + 1;/* endIfGe*/    end
         603 : begin step <= 5043; /* start */ end
         604 : begin if (intermediateValue >= 0) step <=   5097; else step = step + 1;/* endIfGe*/    end
         605 : begin step <= 5084; /* start */ end
         606 : begin if (intermediateValue >= 0) step <=   5138; else step = step + 1;/* endIfGe*/    end
         607 : begin step <= 5125; /* start */ end
         608 : begin if (intermediateValue >= 0) step <=   5179; else step = step + 1;/* endIfGe*/    end
         609 : begin step <= 5166; /* start */ end
         610 : begin if (intermediateValue >= 0) step <=   5220; else step = step + 1;/* endIfGe*/    end
         611 : begin step <= 5207; /* start */ end
         612 : begin if (intermediateValue >= 0) step <=   5261; else step = step + 1;/* endIfGe*/    end
         613 : begin step <= 5248; /* start */ end
         614 : begin if (intermediateValue >= 0) step <=   5302; else step = step + 1;/* endIfGe*/    end
         615 : begin step <= 5289; /* start */ end
         616 : begin if (intermediateValue >= 0) step <=   5343; else step = step + 1;/* endIfGe*/    end
         617 : begin step <= 5330; /* start */ end
         618 : begin if (intermediateValue >= 0) step <=   5384; else step = step + 1;/* endIfGe*/    end
         619 : begin step <= 5371; /* start */ end
         620 : begin memory[196+memory[420]/*mergeRightSibling_r*/]/*free[mergeRightSibling_r]*/ <= -1; /* set 2 */ step <= step + 1; end
         621 : begin memory[217+memory[420]/*mergeRightSibling_r*/]/*isLeaf[mergeRightSibling_r]*/ <= -1; /* set 2 */ step <= step + 1; end
         622 : begin memory[5+memory[420]/*mergeRightSibling_r*/]/*current_size[mergeRightSibling_r]*/ <= -1; /* set 2 */ step <= step + 1; end
         623 : begin memory[196+memory[420]/*mergeRightSibling_r*/]/*free[mergeRightSibling_r]*/ <= intermediateValue; /* set 2 */ step <= step + 1; end
         624 : begin memory[419]/*mergeRightSibling_pk*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         625 : begin intermediateValue <= memory[419]/*mergeRightSibling_pk*/; /* get 1 */ step <= step + 1; end
         626 : begin if (intermediateValue <  0) step <=   5458; else step = step + 1;/* endIfLt*/    end
         627 : begin if (intermediateValue == 0) step <=   5489; else step = step + 1;/* endIfEq*/    end
         628 : begin step <= 5476; /* start */ end
         629 : begin memory[423] <= 1; /* clear 1 */ step <= step + 1; end
         630 : begin step <= 3621; /* start */ end
         631 : begin intermediateValue <= memory[397]/*merge_Key*/; /* get 1 */ step <= step + 1; end
         632 : begin if (intermediateValue >= 0) step <=   5524; else step = step + 1;/* endIfGe*/    end
         633 : begin if (intermediateValue >  0) step <=   5518; else step = step + 1;/* endIfGt*/    end
         634 : begin step <=   5524; /* end */ end
         635 : begin step <= 5508; /* start */ end
         636 : begin intermediateValue <= memory[409]/*merge_loop*/; /* get 1 */ step <= step + 1; end
         637 : begin memory[409]/*merge_loop*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         638 : begin if (intermediateValue >= 0) step <=   5537; else step = step + 1;/* endIfGe*/    end
         639 : begin step <= 3602; /* start */ end
         640 : begin step <=   5869; /* end */ end
         641 : begin if (intermediateValue == 0) step <=   5857; else step = step + 1;/* endIfEq*/    end
         642 : begin memory[445]/*splitBranch_node*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         643 : begin memory[446]/*splitBranch_parent*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         644 : begin memory[443]/*splitBranch_index*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         645 : begin memory[444]/*splitBranch_l*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         646 : begin intermediateValue <= memory[444]/*splitBranch_l*/; /* get 1 */ step <= step + 1; end
         647 : begin if (intermediateValue >  0) step <=   5565; else step = step + 1;/* endIfGt*/    end
         648 : begin intermediateValue <= memory[196+memory[444]/*splitBranch_l*/]/*free[splitBranch_l]*/; /* get 2 */ step <= step + 1; end
         649 : begin memory[196+memory[444]/*splitBranch_l*/]/*free[splitBranch_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         650 : begin memory[217+memory[444]/*splitBranch_l*/]/*isLeaf[splitBranch_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         651 : begin memory[5+memory[444]/*splitBranch_l*/]/*current_size[splitBranch_l]*/ <= 0; /* set 2 */ step <= step + 1; end
         652 : begin intermediateValue <= memory[445]/*splitBranch_node*/; /* get 1 */ step <= step + 1; end
         653 : begin if (intermediateValue >= 0) step <=   5617; else step = step + 1;/* endIfGe*/    end
         654 : begin step <= 5604; /* start */ end
         655 : begin if (intermediateValue >= 0) step <=   5655; else step = step + 1;/* endIfGe*/    end
         656 : begin step <= 5642; /* start */ end
         657 : begin if (intermediateValue >= 0) step <=   5693; else step = step + 1;/* endIfGe*/    end
         658 : begin step <= 5680; /* start */ end
         659 : begin if (intermediateValue >= 0) step <=   5731; else step = step + 1;/* endIfGe*/    end
         660 : begin step <= 5718; /* start */ end
         661 : begin if (intermediateValue >= 0) step <=   5769; else step = step + 1;/* endIfGe*/    end
         662 : begin step <= 5756; /* start */ end
         663 : begin memory[447]/*splitBranch_rk*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         664 : begin intermediateValue <= memory[446]/*splitBranch_parent*/; /* get 1 */ step <= step + 1; end
         665 : begin intermediateValue <= memory[447]/*splitBranch_rk*/; /* get 1 */ step <= step + 1; end
         666 : begin intermediateValue <= memory[443]/*splitBranch_index*/; /* get 1 */ step <= step + 1; end
         667 : begin if (intermediateValue == 0) step <=   5817; else step = step + 1;/* endIfEq*/    end
         668 : begin step <= 5804; /* start */ end
         669 : begin if (intermediateValue >= 0) step <=   5851; else step = step + 1;/* endIfGe*/    end
         670 : begin if (intermediateValue >  0) step <=   5845; else step = step + 1;/* endIfGt*/    end
         671 : begin step <=   5851; /* end */ end
         672 : begin step <= 5835; /* start */ end
         673 : begin if (intermediateValue >  0) step <=   5861; else step = step + 1;/* endIfGt*/    end
         674 : begin intermediateValue <= memory[434]/*put_loop*/; /* get 1 */ step <= step + 1; end
         675 : begin memory[434]/*put_loop*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         676 : begin if (intermediateValue >  0) step <=   5868; else step = step + 1;/* endIfGt*/    end
         677 : begin step <= 1410; /* start */ end

        default: stopped <= 1;
      endcase
      steps    <= steps + 1;
    end // Execute
  end // Always
endmodule
