//-----------------------------------------------------------------------------
// Generic cpu
// Philip R Brenan at appaapps dot com, Appa Apps Ltd Inc., 2025-01-07
//------------------------------------------------------------------------------
`timescale 10ps/1ps
(* keep_hierarchy = "yes" *)
module put(reset, stop, clock, Key, Data, data, found);                    // Database on a chip
  input                      reset;                                             // Restart the program run sequence when this goes high
  input                      clock;                                             // Program counter clock
  input [16-1:0]  Key;                                             // Input key
  input [16-1:0] Data;                                             // Input data
  output                      stop;                                             // Program has stopped when this goes high
  output[bitsPerInteger-1:0]  data;                                             // Output data
  output                     found;                                             // Whether the key was found on put, find delete


  always @ (posedge clock) begin                                                // Execute next step in program
    if (reset) begin                                                            // Reset
      step     <= 0;
      steps    <= 0;
      stopped  <= 0;
    end
    else begin                                                                  // Run
        steps <= steps + 1;
        case(step)
           0: begin intermediateValue = memory[285]; /* get 1 */ end
           1: begin memory[111] = 0; /*set 1 */ end
           2: begin intermediateValue = memory[284]; /* get 1 */ end
           3: begin memory[110] = 0; /*set 1 */ end
           4: begin intermediateValue = memory[111]; /* get 1 */ end
           5: begin memory[113] = 0; /*set 1 */ end
           6: begin intermediateValue = memory[145]; /* get 2 */ end
           7: begin memory[288] = 0; /*set 1 */ end
           8: begin intermediateValue = memory[288]; /* get 1 */ end
           9: begin if (intermediateValue == 0) step =   end.instruction-1; end
          10: begin memory[348] = 0; /*set 1 */ end
          11: begin intermediateValue = memory[113]; /* get 1 */ end
          12: begin memory[294] = 0; /*set 1 */ end
          13: begin memory[292] = 0; /*set 1 */ end
          14: begin memory[293] = 0; /*set 1 */ end
          15: begin intermediateValue = memory[5]; /* get 2 */ end
          16: begin memory[344] = 0; /*set 1 */ end
          17: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
          18: begin if (intermediateValue >= 0) step =   end.instruction-1; end
          19: begin intermediateValue = memory[294]; < memory[166]; ? -1 : memory[294]; == memory[166]; ?  0 : +1; /* compare 2 */ end
          20: begin if (intermediateValue != 0) step =   end.instruction-1; end
          21: begin memory[292] = 1; /*set 1 */ end
          22: begin intermediateValue = memory[166]; /* get 3 */ end
          23: begin memory[294] = 0; /*set 1 */ end
          24: begin intermediateValue = memory[25]; /* get 3 */ end
          25: begin memory[289] = 0; /*set 1 */ end
          26: begin step =   end.instruction-1; end
          27: begin intermediateValue = memory[293]; /* get 1 */ end
          28: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
          29: begin memory[293] = 0; /*set 1 */ end
          30: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
          31: begin if (intermediateValue >= 0) step =   end.instruction-1; end
          32: begin step = start.instruction-1; end
          33: begin intermediateValue = memory[287]; /* get 1 */ end
          34: begin memory[118] = 0; /*set 1 */ end
          35: begin intermediateValue = memory[292]; /* get 1 */ end
          36: begin memory[108] = 0; /*set 1 */ end
          37: begin intermediateValue = memory[293]; /* get 1 */ end
          38: begin memory[112] = 0; /*set 1 */ end
          39: begin intermediateValue = memory[294]; /* get 1 */ end
          40: begin memory[117] = 0; /*set 1 */ end
          41: begin intermediateValue = memory[289]; /* get 1 */ end
          42: begin memory[107] = 0; /*set 1 */ end
          43: begin step =   end.instruction-1; end
          44: begin intermediateValue = memory[287]; /* get 1 */ end
          45: begin memory[283] = 0; /*set 1 */ end
          46: begin memory[114] = 0; /* clear 1 */ end
          47: begin intermediateValue = memory[283]; /* get 1 */ end
          48: begin memory[348] = 0; /*set 1 */ end
          49: begin intermediateValue = memory[113]; /* get 1 */ end
          50: begin memory[294] = 0; /*set 1 */ end
          51: begin memory[292] = 0; /*set 1 */ end
          52: begin memory[293] = 0; /*set 1 */ end
          53: begin intermediateValue = memory[5]; /* get 2 */ end
          54: begin memory[344] = 0; /*set 1 */ end
          55: begin intermediateValue = memory[344]; /* get 1 */ end
          56: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
          57: begin memory[344] = 0; /*set 1 */ end
          58: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
          59: begin if (intermediateValue >= 0) step =   end.instruction-1; end
          60: begin intermediateValue = memory[294]; < memory[166]; ? -1 : memory[294]; == memory[166]; ?  0 : +1; /* compare 2 */ end
          61: begin if (intermediateValue >  0) step =   end.instruction-1; end
          62: begin memory[292] = 1; /*set 1 */ end
          63: begin intermediateValue = memory[166]; /* get 3 */ end
          64: begin memory[294] = 0; /*set 1 */ end
          65: begin intermediateValue = memory[25]; /* get 3 */ end
          66: begin memory[289] = 0; /*set 1 */ end
          67: begin step =   end.instruction-1; end
          68: begin intermediateValue = memory[293]; /* get 1 */ end
          69: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
          70: begin memory[293] = 0; /*set 1 */ end
          71: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
          72: begin if (intermediateValue >= 0) step =   end.instruction-1; end
          73: begin step = start.instruction-1; end
          74: begin intermediateValue = memory[166]; /* get 3 */ end
          75: begin memory[294] = 0; /*set 1 */ end
          76: begin intermediateValue = memory[25]; /* get 3 */ end
          77: begin memory[289] = 0; /*set 1 */ end
          78: begin intermediateValue = memory[289]; /* get 1 */ end
          79: begin memory[4] = 0; /*set 1 */ end
          80: begin intermediateValue = memory[4]; /* get 1 */ end
          81: begin memory[142] = 0; /*set 1 */ end
          82: begin intermediateValue = memory[145]; /* get 2 */ end
          83: begin memory[142] = 0; /*set 1 */ end
          84: begin intermediateValue = memory[142]; /* get 1 */ end
          85: begin if (intermediateValue == 0) step =   end.instruction-1; end
          86: begin intermediateValue = memory[4]; /* get 1 */ end
          87: begin memory[348] = 0; /*set 1 */ end
          88: begin intermediateValue = memory[113]; /* get 1 */ end
          89: begin memory[294] = 0; /*set 1 */ end
          90: begin memory[292] = 0; /*set 1 */ end
          91: begin memory[293] = 0; /*set 1 */ end
          92: begin intermediateValue = memory[5]; /* get 2 */ end
          93: begin memory[344] = 0; /*set 1 */ end
          94: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
          95: begin if (intermediateValue >= 0) step =   end.instruction-1; end
          96: begin intermediateValue = memory[294]; < memory[166]; ? -1 : memory[294]; == memory[166]; ?  0 : +1; /* compare 2 */ end
          97: begin if (intermediateValue != 0) step =   end.instruction-1; end
          98: begin memory[292] = 1; /*set 1 */ end
          99: begin intermediateValue = memory[166]; /* get 3 */ end
         100: begin memory[294] = 0; /*set 1 */ end
         101: begin intermediateValue = memory[25]; /* get 3 */ end
         102: begin memory[289] = 0; /*set 1 */ end
         103: begin step =   end.instruction-1; end
         104: begin intermediateValue = memory[293]; /* get 1 */ end
         105: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         106: begin memory[293] = 0; /*set 1 */ end
         107: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
         108: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         109: begin step = start.instruction-1; end
         110: begin intermediateValue = memory[4]; /* get 1 */ end
         111: begin memory[115] = 0; /*set 1 */ end
         112: begin intermediateValue = memory[115]; /* get 1 */ end
         113: begin memory[118] = 0; /*set 1 */ end
         114: begin intermediateValue = memory[292]; /* get 1 */ end
         115: begin memory[108] = 0; /*set 1 */ end
         116: begin intermediateValue = memory[293]; /* get 1 */ end
         117: begin memory[112] = 0; /*set 1 */ end
         118: begin intermediateValue = memory[294]; /* get 1 */ end
         119: begin memory[117] = 0; /*set 1 */ end
         120: begin intermediateValue = memory[289]; /* get 1 */ end
         121: begin memory[107] = 0; /*set 1 */ end
         122: begin step =   end.instruction-1; end
         123: begin intermediateValue = memory[4]; /* get 1 */ end
         124: begin memory[283] = 0; /*set 1 */ end
         125: begin intermediateValue = memory[114]; /* get 1 */ end
         126: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         127: begin memory[114] = 0; /*set 1 */ end
         128: begin intermediateValue = memory[114]; /* get 1 */ end
         129: begin intermediateValue = 9 <  intermediateValue ? -1 : 9 == intermediateValue ?  0 : +1; /* compare 1 */ end
         130: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         131: begin step = start.instruction-1; end
         132: begin $finish("Search did not terminate in a leaf"); end
         133: begin intermediateValue = memory[108]; /* get 1 */ end
         134: begin if (intermediateValue == 0) step =   end.instruction-1; end
         135: begin intermediateValue = memory[118]; /* get 1 */ end
         136: begin memory[348] = 0; /*set 1 */ end
         137: begin intermediateValue = memory[111]; /* get 1 */ end
         138: begin memory[294] = 0; /*set 1 */ end
         139: begin intermediateValue = memory[110]; /* get 1 */ end
         140: begin memory[289] = 0; /*set 1 */ end
         141: begin intermediateValue = memory[112]; /* get 1 */ end
         142: begin memory[293] = 0; /*set 1 */ end
         143: begin intermediateValue = memory[294]; /* get 1 */ end
         144: begin memory[166] = 0; /*set 3 */ end
         145: begin intermediateValue = memory[289]; /* get 1 */ end
         146: begin memory[25] = 0; /*set 3 */ end
         147: begin intermediateValue = memory[293]; < memory[5]; ? -1 : memory[293]; == memory[5]; ?  0 : +1; /* compare 2 */ end
         148: begin if (intermediateValue <  0) step =   end.instruction-1; end
         149: begin intermediateValue = memory[5]; /* get 2 */ end
         150: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         151: begin memory[5] = 0; /*set 2 */ end
         152: begin memory[140] = 1; /*set 1 */ end
         153: begin memory[116] = 0; /*set 1 */ end
         154: begin step =   end.instruction-1; end
         155: begin intermediateValue = memory[118]; /* get 1 */ end
         156: begin memory[144] = 0; /*set 1 */ end
         157: begin intermediateValue = memory[144]; /* get 1 */ end
         158: begin memory[246] = 0; /*set 1 */ end
         159: begin intermediateValue = memory[5]; /* get 2 */ end
         160: begin memory[246] = 0; /*set 1 */ end
         161: begin intermediateValue = memory[246]; /* get 1 */ end
         162: begin intermediateValue = 2 <  intermediateValue ? -1 : 2 == intermediateValue ?  0 : +1; /* compare 1 */ end
         163: begin intermediateValue = intermediateValue >= 0 ? 1 : 0; /* ge */ end
         164: begin memory[144] = 0; /*set 1 */ end
         165: begin intermediateValue = memory[144]; /* get 1 */ end
         166: begin if (intermediateValue >  0) step =   end.instruction-1; end
         167: begin intermediateValue = memory[118]; /* get 1 */ end
         168: begin memory[348] = 0; /*set 1 */ end
         169: begin intermediateValue = memory[111]; /* get 1 */ end
         170: begin memory[294] = 0; /*set 1 */ end
         171: begin memory[292] = 0; /*set 1 */ end
         172: begin memory[293] = 0; /*set 1 */ end
         173: begin intermediateValue = memory[5]; /* get 2 */ end
         174: begin memory[344] = 0; /*set 1 */ end
         175: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
         176: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         177: begin intermediateValue = memory[294]; < memory[166]; ? -1 : memory[294]; == memory[166]; ?  0 : +1; /* compare 2 */ end
         178: begin if (intermediateValue >  0) step =   end.instruction-1; end
         179: begin memory[292] = 1; /*set 1 */ end
         180: begin intermediateValue = memory[166]; /* get 3 */ end
         181: begin memory[294] = 0; /*set 1 */ end
         182: begin intermediateValue = memory[25]; /* get 3 */ end
         183: begin memory[289] = 0; /*set 1 */ end
         184: begin step =   end.instruction-1; end
         185: begin intermediateValue = memory[293]; /* get 1 */ end
         186: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         187: begin memory[293] = 0; /*set 1 */ end
         188: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
         189: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         190: begin step = start.instruction-1; end
         191: begin intermediateValue = memory[118]; /* get 1 */ end
         192: begin memory[348] = 0; /*set 1 */ end
         193: begin intermediateValue = memory[111]; /* get 1 */ end
         194: begin memory[294] = 0; /*set 1 */ end
         195: begin intermediateValue = memory[110]; /* get 1 */ end
         196: begin memory[289] = 0; /*set 1 */ end
         197: begin intermediateValue = memory[293]; /* get 1 */ end
         198: begin memory[340] = 0; /*set 1 */ end
         199: begin intermediateValue = memory[5]; /* get 2 */ end
         200: begin memory[339] = 0; /*set 1 */ end
         201: begin intermediateValue = memory[339]; /* get 1 */ end
         202: begin memory[338] = 0; /*set 1 */ end
         203: begin intermediateValue = memory[338]; /* get 1 */ end
         204: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
         205: begin memory[338] = 0; /*set 1 */ end
         206: begin intermediateValue = memory[339]; < memory[340]; ? -1 : memory[339]; == memory[340]; ?  0 : +1; /* compare 2 */ end
         207: begin if (intermediateValue == 0) step =   end.instruction-1; end
         208: begin intermediateValue = memory[166]; /* get 3 */ end
         209: begin memory[166] = 0; /*set 3 */ end
         210: begin intermediateValue = memory[25]; /* get 3 */ end
         211: begin memory[25] = 0; /*set 3 */ end
         212: begin intermediateValue = memory[339]; /* get 1 */ end
         213: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
         214: begin memory[339] = 0; /*set 1 */ end
         215: begin intermediateValue = memory[338]; /* get 1 */ end
         216: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
         217: begin memory[338] = 0; /*set 1 */ end
         218: begin step = start.instruction-1; end
         219: begin intermediateValue = memory[294]; /* get 1 */ end
         220: begin memory[166] = 0; /*set 3 */ end
         221: begin intermediateValue = memory[289]; /* get 1 */ end
         222: begin memory[25] = 0; /*set 3 */ end
         223: begin intermediateValue = memory[5]; /* get 2 */ end
         224: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         225: begin memory[5] = 0; /*set 2 */ end
         226: begin memory[140] = 1; /*set 1 */ end
         227: begin memory[116] = 0; /*set 1 */ end
         228: begin step =   end.instruction-1; end
         229: begin memory[140] = 0; /*set 1 */ end
         230: begin memory[116] = 0; /*set 1 */ end
         231: begin intermediateValue = memory[140]; /* get 1 */ end
         232: begin if (intermediateValue >  0) step =   end.instruction-1; end
         233: begin memory[144] = 0; /* clear 1 */ end
         234: begin intermediateValue = memory[144]; /* get 1 */ end
         235: begin memory[142] = 0; /*set 1 */ end
         236: begin intermediateValue = memory[145]; /* get 2 */ end
         237: begin memory[142] = 0; /*set 1 */ end
         238: begin intermediateValue = memory[142]; /* get 1 */ end
         239: begin if (intermediateValue == 0) step =   end.instruction-1; end
         240: begin intermediateValue = memory[144]; /* get 1 */ end
         241: begin memory[246] = 0; /*set 1 */ end
         242: begin intermediateValue = memory[5]; /* get 2 */ end
         243: begin memory[246] = 0; /*set 1 */ end
         244: begin intermediateValue = memory[246]; /* get 1 */ end
         245: begin intermediateValue = 2 <  intermediateValue ? -1 : 2 == intermediateValue ?  0 : +1; /* compare 1 */ end
         246: begin intermediateValue = intermediateValue >= 0 ? 1 : 0; /* ge */ end
         247: begin memory[144] = 0; /*set 1 */ end
         248: begin if (intermediateValue >  0) step =   end.instruction-1; end
         249: begin intermediateValue = memory[144]; /* get 1 */ end
         250: begin memory[3] = 0; /*set 1 */ end
         251: begin intermediateValue = memory[5]; /* get 2 */ end
         252: begin memory[3] = 0; /*set 1 */ end
         253: begin intermediateValue = memory[3]; /* get 1 */ end
         254: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
         255: begin memory[3] = 0; /*set 1 */ end
         256: begin intermediateValue = memory[3]; /* get 1 */ end
         257: begin intermediateValue = 3 <  intermediateValue ? -1 : 3 == intermediateValue ?  0 : +1; /* compare 1 */ end
         258: begin intermediateValue = intermediateValue >= 0 ? 1 : 0; /* ge */ end
         259: begin memory[144] = 0; /*set 1 */ end
         260: begin intermediateValue = memory[144]; /* get 1 */ end
         261: begin memory[143] = 0; /*set 1 */ end
         262: begin intermediateValue = memory[143]; /* get 1 */ end
         263: begin if (intermediateValue == 0) step =   end.instruction-1; end
         264: begin intermediateValue = memory[145]; /* get 2 */ end
         265: begin memory[288] = 0; /*set 1 */ end
         266: begin intermediateValue = memory[288]; /* get 1 */ end
         267: begin if (intermediateValue == 0) step =   end.instruction-1; end
         268: begin intermediateValue = memory[119]; /* get 1 */ end
         269: begin memory[314] = 0; /*set 1 */ end
         270: begin intermediateValue = memory[314]; /* get 1 */ end
         271: begin if (intermediateValue >  0) step =   end.instruction-1; end
         272: begin $finish("No more memory available"); end
         273: begin intermediateValue = memory[120]; /* get 2 */ end
         274: begin memory[119] = 0; /*set 1 */ end
         275: begin memory[120] = 0; /*set 2 */ end
         276: begin memory[145] = 0; /*set 2 */ end
         277: begin memory[5] = 0; /*set 2 */ end
         278: begin memory[166] = 0; /* clear 2 */ end
         279: begin memory[167] = 0; /* clear 2 */ end
         280: begin memory[168] = 0; /* clear 2 */ end
         281: begin memory[169] = 0; /* clear 2 */ end
         282: begin memory[25] = 0; /* clear 2 */ end
         283: begin memory[26] = 0; /* clear 2 */ end
         284: begin memory[27] = 0; /* clear 2 */ end
         285: begin memory[28] = 0; /* clear 2 */ end
         286: begin intermediateValue = memory[314]; /* get 1 */ end
         287: begin memory[291] = 0; /*set 1 */ end
         288: begin memory[145] = 1; /*set 2 */ end
         289: begin intermediateValue = memory[119]; /* get 1 */ end
         290: begin memory[315] = 0; /*set 1 */ end
         291: begin intermediateValue = memory[315]; /* get 1 */ end
         292: begin if (intermediateValue >  0) step =   end.instruction-1; end
         293: begin $finish("No more memory available"); end
         294: begin intermediateValue = memory[120]; /* get 2 */ end
         295: begin memory[119] = 0; /*set 1 */ end
         296: begin memory[120] = 0; /*set 2 */ end
         297: begin memory[145] = 0; /*set 2 */ end
         298: begin memory[5] = 0; /*set 2 */ end
         299: begin memory[166] = 0; /* clear 2 */ end
         300: begin memory[167] = 0; /* clear 2 */ end
         301: begin memory[168] = 0; /* clear 2 */ end
         302: begin memory[169] = 0; /* clear 2 */ end
         303: begin memory[25] = 0; /* clear 2 */ end
         304: begin memory[26] = 0; /* clear 2 */ end
         305: begin memory[27] = 0; /* clear 2 */ end
         306: begin memory[28] = 0; /* clear 2 */ end
         307: begin intermediateValue = memory[315]; /* get 1 */ end
         308: begin memory[291] = 0; /*set 1 */ end
         309: begin memory[145] = 1; /*set 2 */ end
         310: begin intermediateValue = memory[287]; /* get 1 */ end
         311: begin memory[348] = 0; /*set 1 */ end
         312: begin memory[293] = 0; /* clear 1 */ end
         313: begin intermediateValue = memory[166]; /* get 3 */ end
         314: begin memory[294] = 0; /*set 1 */ end
         315: begin intermediateValue = memory[25]; /* get 3 */ end
         316: begin memory[289] = 0; /*set 1 */ end
         317: begin intermediateValue = memory[5]; /* get 2 */ end
         318: begin memory[347] = 0; /*set 1 */ end
         319: begin memory[345] = 0; /*set 1 */ end
         320: begin memory[346] = 1; /*set 1 */ end
         321: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
         322: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         323: begin intermediateValue = memory[166]; /* get 3 */ end
         324: begin memory[166] = 0; /*set 3 */ end
         325: begin intermediateValue = memory[25]; /* get 3 */ end
         326: begin memory[25] = 0; /*set 3 */ end
         327: begin intermediateValue = memory[345]; /* get 1 */ end
         328: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         329: begin memory[345] = 0; /*set 1 */ end
         330: begin intermediateValue = memory[346]; /* get 1 */ end
         331: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         332: begin memory[346] = 0; /*set 1 */ end
         333: begin step = start.instruction-1; end
         334: begin intermediateValue = memory[5]; /* get 2 */ end
         335: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
         336: begin memory[5] = 0; /*set 2 */ end
         337: begin intermediateValue = memory[314]; /* get 1 */ end
         338: begin memory[348] = 0; /*set 1 */ end
         339: begin intermediateValue = memory[5]; /* get 2 */ end
         340: begin memory[293] = 0; /*set 1 */ end
         341: begin intermediateValue = memory[294]; /* get 1 */ end
         342: begin memory[166] = 0; /*set 3 */ end
         343: begin intermediateValue = memory[289]; /* get 1 */ end
         344: begin memory[25] = 0; /*set 3 */ end
         345: begin intermediateValue = memory[5]; /* get 2 */ end
         346: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         347: begin memory[5] = 0; /*set 2 */ end
         348: begin intermediateValue = memory[287]; /* get 1 */ end
         349: begin memory[348] = 0; /*set 1 */ end
         350: begin memory[293] = 0; /* clear 1 */ end
         351: begin intermediateValue = memory[166]; /* get 3 */ end
         352: begin memory[294] = 0; /*set 1 */ end
         353: begin intermediateValue = memory[25]; /* get 3 */ end
         354: begin memory[289] = 0; /*set 1 */ end
         355: begin intermediateValue = memory[5]; /* get 2 */ end
         356: begin memory[347] = 0; /*set 1 */ end
         357: begin memory[345] = 0; /*set 1 */ end
         358: begin memory[346] = 1; /*set 1 */ end
         359: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
         360: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         361: begin intermediateValue = memory[166]; /* get 3 */ end
         362: begin memory[166] = 0; /*set 3 */ end
         363: begin intermediateValue = memory[25]; /* get 3 */ end
         364: begin memory[25] = 0; /*set 3 */ end
         365: begin intermediateValue = memory[345]; /* get 1 */ end
         366: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         367: begin memory[345] = 0; /*set 1 */ end
         368: begin intermediateValue = memory[346]; /* get 1 */ end
         369: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         370: begin memory[346] = 0; /*set 1 */ end
         371: begin step = start.instruction-1; end
         372: begin intermediateValue = memory[5]; /* get 2 */ end
         373: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
         374: begin memory[5] = 0; /*set 2 */ end
         375: begin intermediateValue = memory[315]; /* get 1 */ end
         376: begin memory[348] = 0; /*set 1 */ end
         377: begin intermediateValue = memory[5]; /* get 2 */ end
         378: begin memory[293] = 0; /*set 1 */ end
         379: begin intermediateValue = memory[294]; /* get 1 */ end
         380: begin memory[166] = 0; /*set 3 */ end
         381: begin intermediateValue = memory[289]; /* get 1 */ end
         382: begin memory[25] = 0; /*set 3 */ end
         383: begin intermediateValue = memory[5]; /* get 2 */ end
         384: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         385: begin memory[5] = 0; /*set 2 */ end
         386: begin memory[293] = 0; /*set 1 */ end
         387: begin intermediateValue = memory[166]; /* get 3 */ end
         388: begin memory[294] = 0; /*set 1 */ end
         389: begin intermediateValue = memory[25]; /* get 3 */ end
         390: begin memory[289] = 0; /*set 1 */ end
         391: begin intermediateValue = memory[294]; /* get 1 */ end
         392: begin memory[310] = 0; /*set 1 */ end
         393: begin intermediateValue = memory[314]; /* get 1 */ end
         394: begin memory[348] = 0; /*set 1 */ end
         395: begin intermediateValue = memory[5]; /* get 2 */ end
         396: begin memory[293] = 0; /*set 1 */ end
         397: begin intermediateValue = memory[293]; /* get 1 */ end
         398: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
         399: begin memory[293] = 0; /*set 1 */ end
         400: begin intermediateValue = memory[166]; /* get 3 */ end
         401: begin memory[294] = 0; /*set 1 */ end
         402: begin intermediateValue = memory[25]; /* get 3 */ end
         403: begin memory[289] = 0; /*set 1 */ end
         404: begin intermediateValue = memory[294]; /* get 1 */ end
         405: begin memory[313] = 0; /*set 1 */ end
         406: begin intermediateValue = memory[313]; /* get 1 */ end
         407: begin memory[312] = 0; /*set 1 */ end
         408: begin intermediateValue  = memory[310]; + memory[312];; /* add2 */ end
         409: begin memory[312] = 0; /*set 1 */ end
         410: begin intermediateValue = memory[312]; /* get 1 */ end
         411: begin intermediateValue = intermediateValue >> 1; /* shift right */ end
         412: begin memory[312] = 0; /*set 1 */ end
         413: begin memory[145] = 0; /*set 2 */ end
         414: begin intermediateValue = memory[287]; /* get 1 */ end
         415: begin memory[348] = 0; /*set 1 */ end
         416: begin memory[5] = 0; /*set 2 */ end
         417: begin intermediateValue = memory[312]; /* get 1 */ end
         418: begin memory[294] = 0; /*set 1 */ end
         419: begin intermediateValue = memory[314]; /* get 1 */ end
         420: begin memory[289] = 0; /*set 1 */ end
         421: begin intermediateValue = memory[5]; /* get 2 */ end
         422: begin memory[293] = 0; /*set 1 */ end
         423: begin intermediateValue = memory[294]; /* get 1 */ end
         424: begin memory[166] = 0; /*set 3 */ end
         425: begin intermediateValue = memory[289]; /* get 1 */ end
         426: begin memory[25] = 0; /*set 3 */ end
         427: begin intermediateValue = memory[5]; /* get 2 */ end
         428: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         429: begin memory[5] = 0; /*set 2 */ end
         430: begin intermediateValue = memory[287]; /* get 1 */ end
         431: begin memory[294] = 0; /*set 1 */ end
         432: begin intermediateValue = memory[315]; /* get 1 */ end
         433: begin memory[289] = 0; /*set 1 */ end
         434: begin intermediateValue = memory[5]; /* get 2 */ end
         435: begin memory[293] = 0; /*set 1 */ end
         436: begin intermediateValue = memory[294]; /* get 1 */ end
         437: begin memory[166] = 0; /*set 3 */ end
         438: begin intermediateValue = memory[289]; /* get 1 */ end
         439: begin memory[25] = 0; /*set 3 */ end
         440: begin intermediateValue = memory[5]; /* get 2 */ end
         441: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         442: begin memory[5] = 0; /*set 2 */ end
         443: begin intermediateValue = memory[288]; /* get 1 */ end
         444: begin if (intermediateValue >  0) step =   end.instruction-1; end
         445: begin intermediateValue = memory[119]; /* get 1 */ end
         446: begin memory[300] = 0; /*set 1 */ end
         447: begin intermediateValue = memory[300]; /* get 1 */ end
         448: begin if (intermediateValue >  0) step =   end.instruction-1; end
         449: begin $finish("No more memory available"); end
         450: begin intermediateValue = memory[120]; /* get 2 */ end
         451: begin memory[119] = 0; /*set 1 */ end
         452: begin memory[120] = 0; /*set 2 */ end
         453: begin memory[145] = 0; /*set 2 */ end
         454: begin memory[5] = 0; /*set 2 */ end
         455: begin memory[166] = 0; /* clear 2 */ end
         456: begin memory[167] = 0; /* clear 2 */ end
         457: begin memory[168] = 0; /* clear 2 */ end
         458: begin memory[169] = 0; /* clear 2 */ end
         459: begin memory[25] = 0; /* clear 2 */ end
         460: begin memory[26] = 0; /* clear 2 */ end
         461: begin memory[27] = 0; /* clear 2 */ end
         462: begin memory[28] = 0; /* clear 2 */ end
         463: begin intermediateValue = memory[300]; /* get 1 */ end
         464: begin memory[290] = 0; /*set 1 */ end
         465: begin memory[145] = 0; /*set 2 */ end
         466: begin intermediateValue = memory[119]; /* get 1 */ end
         467: begin memory[302] = 0; /*set 1 */ end
         468: begin intermediateValue = memory[302]; /* get 1 */ end
         469: begin if (intermediateValue >  0) step =   end.instruction-1; end
         470: begin $finish("No more memory available"); end
         471: begin intermediateValue = memory[120]; /* get 2 */ end
         472: begin memory[119] = 0; /*set 1 */ end
         473: begin memory[120] = 0; /*set 2 */ end
         474: begin memory[145] = 0; /*set 2 */ end
         475: begin memory[5] = 0; /*set 2 */ end
         476: begin memory[166] = 0; /* clear 2 */ end
         477: begin memory[167] = 0; /* clear 2 */ end
         478: begin memory[168] = 0; /* clear 2 */ end
         479: begin memory[169] = 0; /* clear 2 */ end
         480: begin memory[25] = 0; /* clear 2 */ end
         481: begin memory[26] = 0; /* clear 2 */ end
         482: begin memory[27] = 0; /* clear 2 */ end
         483: begin memory[28] = 0; /* clear 2 */ end
         484: begin intermediateValue = memory[302]; /* get 1 */ end
         485: begin memory[290] = 0; /*set 1 */ end
         486: begin memory[145] = 0; /*set 2 */ end
         487: begin intermediateValue = memory[287]; /* get 1 */ end
         488: begin memory[348] = 0; /*set 1 */ end
         489: begin memory[293] = 0; /* clear 1 */ end
         490: begin intermediateValue = memory[166]; /* get 3 */ end
         491: begin memory[294] = 0; /*set 1 */ end
         492: begin intermediateValue = memory[25]; /* get 3 */ end
         493: begin memory[289] = 0; /*set 1 */ end
         494: begin intermediateValue = memory[5]; /* get 2 */ end
         495: begin memory[347] = 0; /*set 1 */ end
         496: begin memory[345] = 0; /*set 1 */ end
         497: begin memory[346] = 1; /*set 1 */ end
         498: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
         499: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         500: begin intermediateValue = memory[166]; /* get 3 */ end
         501: begin memory[166] = 0; /*set 3 */ end
         502: begin intermediateValue = memory[25]; /* get 3 */ end
         503: begin memory[25] = 0; /*set 3 */ end
         504: begin intermediateValue = memory[345]; /* get 1 */ end
         505: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         506: begin memory[345] = 0; /*set 1 */ end
         507: begin intermediateValue = memory[346]; /* get 1 */ end
         508: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         509: begin memory[346] = 0; /*set 1 */ end
         510: begin step = start.instruction-1; end
         511: begin intermediateValue = memory[5]; /* get 2 */ end
         512: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
         513: begin memory[5] = 0; /*set 2 */ end
         514: begin intermediateValue = memory[300]; /* get 1 */ end
         515: begin memory[348] = 0; /*set 1 */ end
         516: begin intermediateValue = memory[5]; /* get 2 */ end
         517: begin memory[293] = 0; /*set 1 */ end
         518: begin intermediateValue = memory[294]; /* get 1 */ end
         519: begin memory[166] = 0; /*set 3 */ end
         520: begin intermediateValue = memory[289]; /* get 1 */ end
         521: begin memory[25] = 0; /*set 3 */ end
         522: begin intermediateValue = memory[5]; /* get 2 */ end
         523: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         524: begin memory[5] = 0; /*set 2 */ end
         525: begin intermediateValue = memory[287]; /* get 1 */ end
         526: begin memory[348] = 0; /*set 1 */ end
         527: begin memory[293] = 0; /* clear 1 */ end
         528: begin intermediateValue = memory[166]; /* get 3 */ end
         529: begin memory[294] = 0; /*set 1 */ end
         530: begin intermediateValue = memory[25]; /* get 3 */ end
         531: begin memory[289] = 0; /*set 1 */ end
         532: begin intermediateValue = memory[5]; /* get 2 */ end
         533: begin memory[347] = 0; /*set 1 */ end
         534: begin memory[345] = 0; /*set 1 */ end
         535: begin memory[346] = 1; /*set 1 */ end
         536: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
         537: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         538: begin intermediateValue = memory[166]; /* get 3 */ end
         539: begin memory[166] = 0; /*set 3 */ end
         540: begin intermediateValue = memory[25]; /* get 3 */ end
         541: begin memory[25] = 0; /*set 3 */ end
         542: begin intermediateValue = memory[345]; /* get 1 */ end
         543: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         544: begin memory[345] = 0; /*set 1 */ end
         545: begin intermediateValue = memory[346]; /* get 1 */ end
         546: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         547: begin memory[346] = 0; /*set 1 */ end
         548: begin step = start.instruction-1; end
         549: begin intermediateValue = memory[5]; /* get 2 */ end
         550: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
         551: begin memory[5] = 0; /*set 2 */ end
         552: begin intermediateValue = memory[294]; /* get 1 */ end
         553: begin memory[301] = 0; /*set 1 */ end
         554: begin intermediateValue = memory[300]; /* get 1 */ end
         555: begin memory[348] = 0; /*set 1 */ end
         556: begin intermediateValue = memory[287]; /* get 1 */ end
         557: begin memory[294] = 0; /*set 1 */ end
         558: begin intermediateValue = memory[5]; /* get 2 */ end
         559: begin memory[293] = 0; /*set 1 */ end
         560: begin intermediateValue = memory[294]; /* get 1 */ end
         561: begin memory[166] = 0; /*set 3 */ end
         562: begin intermediateValue = memory[289]; /* get 1 */ end
         563: begin memory[25] = 0; /*set 3 */ end
         564: begin intermediateValue = memory[5]; /* get 2 */ end
         565: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         566: begin memory[5] = 0; /*set 2 */ end
         567: begin intermediateValue = memory[287]; /* get 1 */ end
         568: begin memory[348] = 0; /*set 1 */ end
         569: begin memory[293] = 0; /* clear 1 */ end
         570: begin intermediateValue = memory[166]; /* get 3 */ end
         571: begin memory[294] = 0; /*set 1 */ end
         572: begin intermediateValue = memory[25]; /* get 3 */ end
         573: begin memory[289] = 0; /*set 1 */ end
         574: begin intermediateValue = memory[5]; /* get 2 */ end
         575: begin memory[347] = 0; /*set 1 */ end
         576: begin memory[345] = 0; /*set 1 */ end
         577: begin memory[346] = 1; /*set 1 */ end
         578: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
         579: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         580: begin intermediateValue = memory[166]; /* get 3 */ end
         581: begin memory[166] = 0; /*set 3 */ end
         582: begin intermediateValue = memory[25]; /* get 3 */ end
         583: begin memory[25] = 0; /*set 3 */ end
         584: begin intermediateValue = memory[345]; /* get 1 */ end
         585: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         586: begin memory[345] = 0; /*set 1 */ end
         587: begin intermediateValue = memory[346]; /* get 1 */ end
         588: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         589: begin memory[346] = 0; /*set 1 */ end
         590: begin step = start.instruction-1; end
         591: begin intermediateValue = memory[5]; /* get 2 */ end
         592: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
         593: begin memory[5] = 0; /*set 2 */ end
         594: begin intermediateValue = memory[302]; /* get 1 */ end
         595: begin memory[348] = 0; /*set 1 */ end
         596: begin intermediateValue = memory[5]; /* get 2 */ end
         597: begin memory[293] = 0; /*set 1 */ end
         598: begin intermediateValue = memory[294]; /* get 1 */ end
         599: begin memory[166] = 0; /*set 3 */ end
         600: begin intermediateValue = memory[289]; /* get 1 */ end
         601: begin memory[25] = 0; /*set 3 */ end
         602: begin intermediateValue = memory[5]; /* get 2 */ end
         603: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         604: begin memory[5] = 0; /*set 2 */ end
         605: begin intermediateValue = memory[287]; /* get 1 */ end
         606: begin memory[348] = 0; /*set 1 */ end
         607: begin memory[293] = 0; /* clear 1 */ end
         608: begin intermediateValue = memory[166]; /* get 3 */ end
         609: begin memory[294] = 0; /*set 1 */ end
         610: begin intermediateValue = memory[25]; /* get 3 */ end
         611: begin memory[289] = 0; /*set 1 */ end
         612: begin intermediateValue = memory[5]; /* get 2 */ end
         613: begin memory[347] = 0; /*set 1 */ end
         614: begin memory[345] = 0; /*set 1 */ end
         615: begin memory[346] = 1; /*set 1 */ end
         616: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
         617: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         618: begin intermediateValue = memory[166]; /* get 3 */ end
         619: begin memory[166] = 0; /*set 3 */ end
         620: begin intermediateValue = memory[25]; /* get 3 */ end
         621: begin memory[25] = 0; /*set 3 */ end
         622: begin intermediateValue = memory[345]; /* get 1 */ end
         623: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         624: begin memory[345] = 0; /*set 1 */ end
         625: begin intermediateValue = memory[346]; /* get 1 */ end
         626: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         627: begin memory[346] = 0; /*set 1 */ end
         628: begin step = start.instruction-1; end
         629: begin intermediateValue = memory[5]; /* get 2 */ end
         630: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
         631: begin memory[5] = 0; /*set 2 */ end
         632: begin intermediateValue = memory[302]; /* get 1 */ end
         633: begin memory[348] = 0; /*set 1 */ end
         634: begin intermediateValue = memory[287]; /* get 1 */ end
         635: begin memory[294] = 0; /*set 1 */ end
         636: begin intermediateValue = memory[5]; /* get 2 */ end
         637: begin memory[293] = 0; /*set 1 */ end
         638: begin intermediateValue = memory[294]; /* get 1 */ end
         639: begin memory[166] = 0; /*set 3 */ end
         640: begin intermediateValue = memory[289]; /* get 1 */ end
         641: begin memory[25] = 0; /*set 3 */ end
         642: begin intermediateValue = memory[5]; /* get 2 */ end
         643: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         644: begin memory[5] = 0; /*set 2 */ end
         645: begin intermediateValue = memory[287]; /* get 1 */ end
         646: begin memory[348] = 0; /*set 1 */ end
         647: begin memory[5] = 0; /*set 2 */ end
         648: begin intermediateValue = memory[301]; /* get 1 */ end
         649: begin memory[294] = 0; /*set 1 */ end
         650: begin intermediateValue = memory[300]; /* get 1 */ end
         651: begin memory[289] = 0; /*set 1 */ end
         652: begin intermediateValue = memory[5]; /* get 2 */ end
         653: begin memory[293] = 0; /*set 1 */ end
         654: begin intermediateValue = memory[294]; /* get 1 */ end
         655: begin memory[166] = 0; /*set 3 */ end
         656: begin intermediateValue = memory[289]; /* get 1 */ end
         657: begin memory[25] = 0; /*set 3 */ end
         658: begin intermediateValue = memory[5]; /* get 2 */ end
         659: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         660: begin memory[5] = 0; /*set 2 */ end
         661: begin intermediateValue = memory[287]; /* get 1 */ end
         662: begin memory[294] = 0; /*set 1 */ end
         663: begin intermediateValue = memory[302]; /* get 1 */ end
         664: begin memory[289] = 0; /*set 1 */ end
         665: begin intermediateValue = memory[5]; /* get 2 */ end
         666: begin memory[293] = 0; /*set 1 */ end
         667: begin intermediateValue = memory[294]; /* get 1 */ end
         668: begin memory[166] = 0; /*set 3 */ end
         669: begin intermediateValue = memory[289]; /* get 1 */ end
         670: begin memory[25] = 0; /*set 3 */ end
         671: begin intermediateValue = memory[5]; /* get 2 */ end
         672: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         673: begin memory[5] = 0; /*set 2 */ end
         674: begin intermediateValue = memory[111]; /* get 1 */ end
         675: begin memory[113] = 0; /*set 1 */ end
         676: begin intermediateValue = memory[145]; /* get 2 */ end
         677: begin memory[288] = 0; /*set 1 */ end
         678: begin intermediateValue = memory[288]; /* get 1 */ end
         679: begin if (intermediateValue == 0) step =   end.instruction-1; end
         680: begin memory[348] = 0; /*set 1 */ end
         681: begin intermediateValue = memory[113]; /* get 1 */ end
         682: begin memory[294] = 0; /*set 1 */ end
         683: begin memory[292] = 0; /*set 1 */ end
         684: begin memory[293] = 0; /*set 1 */ end
         685: begin intermediateValue = memory[5]; /* get 2 */ end
         686: begin memory[344] = 0; /*set 1 */ end
         687: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
         688: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         689: begin intermediateValue = memory[294]; < memory[166]; ? -1 : memory[294]; == memory[166]; ?  0 : +1; /* compare 2 */ end
         690: begin if (intermediateValue != 0) step =   end.instruction-1; end
         691: begin memory[292] = 1; /*set 1 */ end
         692: begin intermediateValue = memory[166]; /* get 3 */ end
         693: begin memory[294] = 0; /*set 1 */ end
         694: begin intermediateValue = memory[25]; /* get 3 */ end
         695: begin memory[289] = 0; /*set 1 */ end
         696: begin step =   end.instruction-1; end
         697: begin intermediateValue = memory[293]; /* get 1 */ end
         698: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         699: begin memory[293] = 0; /*set 1 */ end
         700: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
         701: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         702: begin step = start.instruction-1; end
         703: begin intermediateValue = memory[287]; /* get 1 */ end
         704: begin memory[118] = 0; /*set 1 */ end
         705: begin intermediateValue = memory[292]; /* get 1 */ end
         706: begin memory[108] = 0; /*set 1 */ end
         707: begin intermediateValue = memory[293]; /* get 1 */ end
         708: begin memory[112] = 0; /*set 1 */ end
         709: begin intermediateValue = memory[294]; /* get 1 */ end
         710: begin memory[117] = 0; /*set 1 */ end
         711: begin intermediateValue = memory[289]; /* get 1 */ end
         712: begin memory[107] = 0; /*set 1 */ end
         713: begin step =   end.instruction-1; end
         714: begin intermediateValue = memory[287]; /* get 1 */ end
         715: begin memory[283] = 0; /*set 1 */ end
         716: begin memory[114] = 0; /* clear 1 */ end
         717: begin intermediateValue = memory[283]; /* get 1 */ end
         718: begin memory[348] = 0; /*set 1 */ end
         719: begin intermediateValue = memory[113]; /* get 1 */ end
         720: begin memory[294] = 0; /*set 1 */ end
         721: begin memory[292] = 0; /*set 1 */ end
         722: begin memory[293] = 0; /*set 1 */ end
         723: begin intermediateValue = memory[5]; /* get 2 */ end
         724: begin memory[344] = 0; /*set 1 */ end
         725: begin intermediateValue = memory[344]; /* get 1 */ end
         726: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
         727: begin memory[344] = 0; /*set 1 */ end
         728: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
         729: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         730: begin intermediateValue = memory[294]; < memory[166]; ? -1 : memory[294]; == memory[166]; ?  0 : +1; /* compare 2 */ end
         731: begin if (intermediateValue >  0) step =   end.instruction-1; end
         732: begin memory[292] = 1; /*set 1 */ end
         733: begin intermediateValue = memory[166]; /* get 3 */ end
         734: begin memory[294] = 0; /*set 1 */ end
         735: begin intermediateValue = memory[25]; /* get 3 */ end
         736: begin memory[289] = 0; /*set 1 */ end
         737: begin step =   end.instruction-1; end
         738: begin intermediateValue = memory[293]; /* get 1 */ end
         739: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         740: begin memory[293] = 0; /*set 1 */ end
         741: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
         742: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         743: begin step = start.instruction-1; end
         744: begin intermediateValue = memory[166]; /* get 3 */ end
         745: begin memory[294] = 0; /*set 1 */ end
         746: begin intermediateValue = memory[25]; /* get 3 */ end
         747: begin memory[289] = 0; /*set 1 */ end
         748: begin intermediateValue = memory[289]; /* get 1 */ end
         749: begin memory[4] = 0; /*set 1 */ end
         750: begin intermediateValue = memory[4]; /* get 1 */ end
         751: begin memory[142] = 0; /*set 1 */ end
         752: begin intermediateValue = memory[145]; /* get 2 */ end
         753: begin memory[142] = 0; /*set 1 */ end
         754: begin intermediateValue = memory[142]; /* get 1 */ end
         755: begin if (intermediateValue == 0) step =   end.instruction-1; end
         756: begin intermediateValue = memory[4]; /* get 1 */ end
         757: begin memory[348] = 0; /*set 1 */ end
         758: begin intermediateValue = memory[113]; /* get 1 */ end
         759: begin memory[294] = 0; /*set 1 */ end
         760: begin memory[292] = 0; /*set 1 */ end
         761: begin memory[293] = 0; /*set 1 */ end
         762: begin intermediateValue = memory[5]; /* get 2 */ end
         763: begin memory[344] = 0; /*set 1 */ end
         764: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
         765: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         766: begin intermediateValue = memory[294]; < memory[166]; ? -1 : memory[294]; == memory[166]; ?  0 : +1; /* compare 2 */ end
         767: begin if (intermediateValue != 0) step =   end.instruction-1; end
         768: begin memory[292] = 1; /*set 1 */ end
         769: begin intermediateValue = memory[166]; /* get 3 */ end
         770: begin memory[294] = 0; /*set 1 */ end
         771: begin intermediateValue = memory[25]; /* get 3 */ end
         772: begin memory[289] = 0; /*set 1 */ end
         773: begin step =   end.instruction-1; end
         774: begin intermediateValue = memory[293]; /* get 1 */ end
         775: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         776: begin memory[293] = 0; /*set 1 */ end
         777: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
         778: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         779: begin step = start.instruction-1; end
         780: begin intermediateValue = memory[4]; /* get 1 */ end
         781: begin memory[115] = 0; /*set 1 */ end
         782: begin intermediateValue = memory[115]; /* get 1 */ end
         783: begin memory[118] = 0; /*set 1 */ end
         784: begin intermediateValue = memory[292]; /* get 1 */ end
         785: begin memory[108] = 0; /*set 1 */ end
         786: begin intermediateValue = memory[293]; /* get 1 */ end
         787: begin memory[112] = 0; /*set 1 */ end
         788: begin intermediateValue = memory[294]; /* get 1 */ end
         789: begin memory[117] = 0; /*set 1 */ end
         790: begin intermediateValue = memory[289]; /* get 1 */ end
         791: begin memory[107] = 0; /*set 1 */ end
         792: begin step =   end.instruction-1; end
         793: begin intermediateValue = memory[4]; /* get 1 */ end
         794: begin memory[283] = 0; /*set 1 */ end
         795: begin intermediateValue = memory[114]; /* get 1 */ end
         796: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         797: begin memory[114] = 0; /*set 1 */ end
         798: begin intermediateValue = memory[114]; /* get 1 */ end
         799: begin intermediateValue = 9 <  intermediateValue ? -1 : 9 == intermediateValue ?  0 : +1; /* compare 1 */ end
         800: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         801: begin step = start.instruction-1; end
         802: begin $finish("Search did not terminate in a leaf"); end
         803: begin intermediateValue = memory[108]; /* get 1 */ end
         804: begin if (intermediateValue == 0) step =   end.instruction-1; end
         805: begin intermediateValue = memory[118]; /* get 1 */ end
         806: begin memory[348] = 0; /*set 1 */ end
         807: begin intermediateValue = memory[111]; /* get 1 */ end
         808: begin memory[294] = 0; /*set 1 */ end
         809: begin intermediateValue = memory[110]; /* get 1 */ end
         810: begin memory[289] = 0; /*set 1 */ end
         811: begin intermediateValue = memory[112]; /* get 1 */ end
         812: begin memory[293] = 0; /*set 1 */ end
         813: begin intermediateValue = memory[294]; /* get 1 */ end
         814: begin memory[166] = 0; /*set 3 */ end
         815: begin intermediateValue = memory[289]; /* get 1 */ end
         816: begin memory[25] = 0; /*set 3 */ end
         817: begin intermediateValue = memory[293]; < memory[5]; ? -1 : memory[293]; == memory[5]; ?  0 : +1; /* compare 2 */ end
         818: begin if (intermediateValue <  0) step =   end.instruction-1; end
         819: begin intermediateValue = memory[5]; /* get 2 */ end
         820: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         821: begin memory[5] = 0; /*set 2 */ end
         822: begin memory[140] = 1; /*set 1 */ end
         823: begin memory[116] = 0; /*set 1 */ end
         824: begin step =   end.instruction-1; end
         825: begin intermediateValue = memory[118]; /* get 1 */ end
         826: begin memory[144] = 0; /*set 1 */ end
         827: begin intermediateValue = memory[144]; /* get 1 */ end
         828: begin memory[246] = 0; /*set 1 */ end
         829: begin intermediateValue = memory[5]; /* get 2 */ end
         830: begin memory[246] = 0; /*set 1 */ end
         831: begin intermediateValue = memory[246]; /* get 1 */ end
         832: begin intermediateValue = 2 <  intermediateValue ? -1 : 2 == intermediateValue ?  0 : +1; /* compare 1 */ end
         833: begin intermediateValue = intermediateValue >= 0 ? 1 : 0; /* ge */ end
         834: begin memory[144] = 0; /*set 1 */ end
         835: begin intermediateValue = memory[144]; /* get 1 */ end
         836: begin if (intermediateValue >  0) step =   end.instruction-1; end
         837: begin intermediateValue = memory[118]; /* get 1 */ end
         838: begin memory[348] = 0; /*set 1 */ end
         839: begin intermediateValue = memory[111]; /* get 1 */ end
         840: begin memory[294] = 0; /*set 1 */ end
         841: begin memory[292] = 0; /*set 1 */ end
         842: begin memory[293] = 0; /*set 1 */ end
         843: begin intermediateValue = memory[5]; /* get 2 */ end
         844: begin memory[344] = 0; /*set 1 */ end
         845: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
         846: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         847: begin intermediateValue = memory[294]; < memory[166]; ? -1 : memory[294]; == memory[166]; ?  0 : +1; /* compare 2 */ end
         848: begin if (intermediateValue >  0) step =   end.instruction-1; end
         849: begin memory[292] = 1; /*set 1 */ end
         850: begin intermediateValue = memory[166]; /* get 3 */ end
         851: begin memory[294] = 0; /*set 1 */ end
         852: begin intermediateValue = memory[25]; /* get 3 */ end
         853: begin memory[289] = 0; /*set 1 */ end
         854: begin step =   end.instruction-1; end
         855: begin intermediateValue = memory[293]; /* get 1 */ end
         856: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         857: begin memory[293] = 0; /*set 1 */ end
         858: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
         859: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         860: begin step = start.instruction-1; end
         861: begin intermediateValue = memory[118]; /* get 1 */ end
         862: begin memory[348] = 0; /*set 1 */ end
         863: begin intermediateValue = memory[111]; /* get 1 */ end
         864: begin memory[294] = 0; /*set 1 */ end
         865: begin intermediateValue = memory[110]; /* get 1 */ end
         866: begin memory[289] = 0; /*set 1 */ end
         867: begin intermediateValue = memory[293]; /* get 1 */ end
         868: begin memory[340] = 0; /*set 1 */ end
         869: begin intermediateValue = memory[5]; /* get 2 */ end
         870: begin memory[339] = 0; /*set 1 */ end
         871: begin intermediateValue = memory[339]; /* get 1 */ end
         872: begin memory[338] = 0; /*set 1 */ end
         873: begin intermediateValue = memory[338]; /* get 1 */ end
         874: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
         875: begin memory[338] = 0; /*set 1 */ end
         876: begin intermediateValue = memory[339]; < memory[340]; ? -1 : memory[339]; == memory[340]; ?  0 : +1; /* compare 2 */ end
         877: begin if (intermediateValue == 0) step =   end.instruction-1; end
         878: begin intermediateValue = memory[166]; /* get 3 */ end
         879: begin memory[166] = 0; /*set 3 */ end
         880: begin intermediateValue = memory[25]; /* get 3 */ end
         881: begin memory[25] = 0; /*set 3 */ end
         882: begin intermediateValue = memory[339]; /* get 1 */ end
         883: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
         884: begin memory[339] = 0; /*set 1 */ end
         885: begin intermediateValue = memory[338]; /* get 1 */ end
         886: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
         887: begin memory[338] = 0; /*set 1 */ end
         888: begin step = start.instruction-1; end
         889: begin intermediateValue = memory[294]; /* get 1 */ end
         890: begin memory[166] = 0; /*set 3 */ end
         891: begin intermediateValue = memory[289]; /* get 1 */ end
         892: begin memory[25] = 0; /*set 3 */ end
         893: begin intermediateValue = memory[5]; /* get 2 */ end
         894: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         895: begin memory[5] = 0; /*set 2 */ end
         896: begin memory[140] = 1; /*set 1 */ end
         897: begin memory[116] = 0; /*set 1 */ end
         898: begin step =   end.instruction-1; end
         899: begin memory[140] = 0; /*set 1 */ end
         900: begin memory[116] = 0; /*set 1 */ end
         901: begin intermediateValue = memory[140]; /* get 1 */ end
         902: begin if (intermediateValue >  0) step =   end.instruction-1; end
         903: begin intermediateValue = memory[287]; /* get 1 */ end
         904: begin memory[283] = 0; /*set 1 */ end
         905: begin memory[286] = 0; /* clear 1 */ end
         906: begin intermediateValue = memory[283]; /* get 1 */ end
         907: begin memory[348] = 0; /*set 1 */ end
         908: begin intermediateValue = memory[285]; /* get 1 */ end
         909: begin memory[294] = 0; /*set 1 */ end
         910: begin memory[292] = 0; /*set 1 */ end
         911: begin memory[293] = 0; /*set 1 */ end
         912: begin intermediateValue = memory[5]; /* get 2 */ end
         913: begin memory[344] = 0; /*set 1 */ end
         914: begin intermediateValue = memory[344]; /* get 1 */ end
         915: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
         916: begin memory[344] = 0; /*set 1 */ end
         917: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
         918: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         919: begin intermediateValue = memory[294]; < memory[166]; ? -1 : memory[294]; == memory[166]; ?  0 : +1; /* compare 2 */ end
         920: begin if (intermediateValue >  0) step =   end.instruction-1; end
         921: begin memory[292] = 1; /*set 1 */ end
         922: begin intermediateValue = memory[166]; /* get 3 */ end
         923: begin memory[294] = 0; /*set 1 */ end
         924: begin intermediateValue = memory[25]; /* get 3 */ end
         925: begin memory[289] = 0; /*set 1 */ end
         926: begin step =   end.instruction-1; end
         927: begin intermediateValue = memory[293]; /* get 1 */ end
         928: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         929: begin memory[293] = 0; /*set 1 */ end
         930: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
         931: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         932: begin step = start.instruction-1; end
         933: begin intermediateValue = memory[166]; /* get 3 */ end
         934: begin memory[294] = 0; /*set 1 */ end
         935: begin intermediateValue = memory[25]; /* get 3 */ end
         936: begin memory[289] = 0; /*set 1 */ end
         937: begin intermediateValue = memory[289]; /* get 1 */ end
         938: begin memory[4] = 0; /*set 1 */ end
         939: begin intermediateValue = memory[4]; /* get 1 */ end
         940: begin memory[142] = 0; /*set 1 */ end
         941: begin intermediateValue = memory[145]; /* get 2 */ end
         942: begin memory[142] = 0; /*set 1 */ end
         943: begin intermediateValue = memory[142]; /* get 1 */ end
         944: begin if (intermediateValue == 0) step =   end.instruction-1; end
         945: begin intermediateValue = memory[4]; /* get 1 */ end
         946: begin memory[308] = 0; /*set 1 */ end
         947: begin intermediateValue = memory[283]; /* get 1 */ end
         948: begin memory[309] = 0; /*set 1 */ end
         949: begin intermediateValue = memory[293]; /* get 1 */ end
         950: begin memory[305] = 0; /*set 1 */ end
         951: begin intermediateValue = memory[119]; /* get 1 */ end
         952: begin memory[307] = 0; /*set 1 */ end
         953: begin intermediateValue = memory[307]; /* get 1 */ end
         954: begin if (intermediateValue >  0) step =   end.instruction-1; end
         955: begin $finish("No more memory available"); end
         956: begin intermediateValue = memory[120]; /* get 2 */ end
         957: begin memory[119] = 0; /*set 1 */ end
         958: begin memory[120] = 0; /*set 2 */ end
         959: begin memory[145] = 0; /*set 2 */ end
         960: begin memory[5] = 0; /*set 2 */ end
         961: begin memory[166] = 0; /* clear 2 */ end
         962: begin memory[167] = 0; /* clear 2 */ end
         963: begin memory[168] = 0; /* clear 2 */ end
         964: begin memory[169] = 0; /* clear 2 */ end
         965: begin memory[25] = 0; /* clear 2 */ end
         966: begin memory[26] = 0; /* clear 2 */ end
         967: begin memory[27] = 0; /* clear 2 */ end
         968: begin memory[28] = 0; /* clear 2 */ end
         969: begin intermediateValue = memory[307]; /* get 1 */ end
         970: begin memory[291] = 0; /*set 1 */ end
         971: begin memory[145] = 1; /*set 2 */ end
         972: begin intermediateValue = memory[308]; /* get 1 */ end
         973: begin memory[348] = 0; /*set 1 */ end
         974: begin memory[293] = 0; /* clear 1 */ end
         975: begin intermediateValue = memory[166]; /* get 3 */ end
         976: begin memory[294] = 0; /*set 1 */ end
         977: begin intermediateValue = memory[25]; /* get 3 */ end
         978: begin memory[289] = 0; /*set 1 */ end
         979: begin intermediateValue = memory[5]; /* get 2 */ end
         980: begin memory[347] = 0; /*set 1 */ end
         981: begin memory[345] = 0; /*set 1 */ end
         982: begin memory[346] = 1; /*set 1 */ end
         983: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
         984: begin if (intermediateValue >= 0) step =   end.instruction-1; end
         985: begin intermediateValue = memory[166]; /* get 3 */ end
         986: begin memory[166] = 0; /*set 3 */ end
         987: begin intermediateValue = memory[25]; /* get 3 */ end
         988: begin memory[25] = 0; /*set 3 */ end
         989: begin intermediateValue = memory[345]; /* get 1 */ end
         990: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         991: begin memory[345] = 0; /*set 1 */ end
         992: begin intermediateValue = memory[346]; /* get 1 */ end
         993: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
         994: begin memory[346] = 0; /*set 1 */ end
         995: begin step = start.instruction-1; end
         996: begin intermediateValue = memory[5]; /* get 2 */ end
         997: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
         998: begin memory[5] = 0; /*set 2 */ end
         999: begin intermediateValue = memory[307]; /* get 1 */ end
        1000: begin memory[348] = 0; /*set 1 */ end
        1001: begin intermediateValue = memory[5]; /* get 2 */ end
        1002: begin memory[293] = 0; /*set 1 */ end
        1003: begin intermediateValue = memory[294]; /* get 1 */ end
        1004: begin memory[166] = 0; /*set 3 */ end
        1005: begin intermediateValue = memory[289]; /* get 1 */ end
        1006: begin memory[25] = 0; /*set 3 */ end
        1007: begin intermediateValue = memory[5]; /* get 2 */ end
        1008: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1009: begin memory[5] = 0; /*set 2 */ end
        1010: begin intermediateValue = memory[308]; /* get 1 */ end
        1011: begin memory[348] = 0; /*set 1 */ end
        1012: begin memory[293] = 0; /*set 1 */ end
        1013: begin intermediateValue = memory[166]; /* get 3 */ end
        1014: begin memory[294] = 0; /*set 1 */ end
        1015: begin intermediateValue = memory[25]; /* get 3 */ end
        1016: begin memory[289] = 0; /*set 1 */ end
        1017: begin intermediateValue = memory[294]; /* get 1 */ end
        1018: begin memory[303] = 0; /*set 1 */ end
        1019: begin intermediateValue = memory[307]; /* get 1 */ end
        1020: begin memory[348] = 0; /*set 1 */ end
        1021: begin intermediateValue = memory[5]; /* get 2 */ end
        1022: begin memory[293] = 0; /*set 1 */ end
        1023: begin intermediateValue = memory[293]; /* get 1 */ end
        1024: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1025: begin memory[293] = 0; /*set 1 */ end
        1026: begin intermediateValue = memory[166]; /* get 3 */ end
        1027: begin memory[294] = 0; /*set 1 */ end
        1028: begin intermediateValue = memory[25]; /* get 3 */ end
        1029: begin memory[289] = 0; /*set 1 */ end
        1030: begin intermediateValue = memory[294]; /* get 1 */ end
        1031: begin memory[306] = 0; /*set 1 */ end
        1032: begin intermediateValue = memory[303]; /* get 1 */ end
        1033: begin memory[304] = 0; /*set 1 */ end
        1034: begin intermediateValue  = memory[306]; + memory[304];; /* add2 */ end
        1035: begin memory[304] = 0; /*set 1 */ end
        1036: begin intermediateValue = memory[304]; /* get 1 */ end
        1037: begin intermediateValue = intermediateValue >> 1; /* shift right */ end
        1038: begin memory[304] = 0; /*set 1 */ end
        1039: begin intermediateValue = memory[309]; /* get 1 */ end
        1040: begin memory[348] = 0; /*set 1 */ end
        1041: begin intermediateValue = memory[304]; /* get 1 */ end
        1042: begin memory[294] = 0; /*set 1 */ end
        1043: begin intermediateValue = memory[307]; /* get 1 */ end
        1044: begin memory[289] = 0; /*set 1 */ end
        1045: begin intermediateValue = memory[305]; /* get 1 */ end
        1046: begin memory[293] = 0; /*set 1 */ end
        1047: begin intermediateValue = memory[293]; /* get 1 */ end
        1048: begin memory[340] = 0; /*set 1 */ end
        1049: begin intermediateValue = memory[5]; /* get 2 */ end
        1050: begin memory[339] = 0; /*set 1 */ end
        1051: begin intermediateValue = memory[339]; /* get 1 */ end
        1052: begin memory[338] = 0; /*set 1 */ end
        1053: begin intermediateValue = memory[338]; /* get 1 */ end
        1054: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1055: begin memory[338] = 0; /*set 1 */ end
        1056: begin intermediateValue = memory[339]; < memory[340]; ? -1 : memory[339]; == memory[340]; ?  0 : +1; /* compare 2 */ end
        1057: begin if (intermediateValue == 0) step =   end.instruction-1; end
        1058: begin intermediateValue = memory[166]; /* get 3 */ end
        1059: begin memory[166] = 0; /*set 3 */ end
        1060: begin intermediateValue = memory[25]; /* get 3 */ end
        1061: begin memory[25] = 0; /*set 3 */ end
        1062: begin intermediateValue = memory[339]; /* get 1 */ end
        1063: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1064: begin memory[339] = 0; /*set 1 */ end
        1065: begin intermediateValue = memory[338]; /* get 1 */ end
        1066: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1067: begin memory[338] = 0; /*set 1 */ end
        1068: begin step = start.instruction-1; end
        1069: begin intermediateValue = memory[294]; /* get 1 */ end
        1070: begin memory[166] = 0; /*set 3 */ end
        1071: begin intermediateValue = memory[289]; /* get 1 */ end
        1072: begin memory[25] = 0; /*set 3 */ end
        1073: begin intermediateValue = memory[5]; /* get 2 */ end
        1074: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1075: begin memory[5] = 0; /*set 2 */ end
        1076: begin intermediateValue = memory[111]; /* get 1 */ end
        1077: begin memory[113] = 0; /*set 1 */ end
        1078: begin intermediateValue = memory[145]; /* get 2 */ end
        1079: begin memory[288] = 0; /*set 1 */ end
        1080: begin intermediateValue = memory[288]; /* get 1 */ end
        1081: begin if (intermediateValue == 0) step =   end.instruction-1; end
        1082: begin memory[348] = 0; /*set 1 */ end
        1083: begin intermediateValue = memory[113]; /* get 1 */ end
        1084: begin memory[294] = 0; /*set 1 */ end
        1085: begin memory[292] = 0; /*set 1 */ end
        1086: begin memory[293] = 0; /*set 1 */ end
        1087: begin intermediateValue = memory[5]; /* get 2 */ end
        1088: begin memory[344] = 0; /*set 1 */ end
        1089: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
        1090: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        1091: begin intermediateValue = memory[294]; < memory[166]; ? -1 : memory[294]; == memory[166]; ?  0 : +1; /* compare 2 */ end
        1092: begin if (intermediateValue != 0) step =   end.instruction-1; end
        1093: begin memory[292] = 1; /*set 1 */ end
        1094: begin intermediateValue = memory[166]; /* get 3 */ end
        1095: begin memory[294] = 0; /*set 1 */ end
        1096: begin intermediateValue = memory[25]; /* get 3 */ end
        1097: begin memory[289] = 0; /*set 1 */ end
        1098: begin step =   end.instruction-1; end
        1099: begin intermediateValue = memory[293]; /* get 1 */ end
        1100: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1101: begin memory[293] = 0; /*set 1 */ end
        1102: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
        1103: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        1104: begin step = start.instruction-1; end
        1105: begin intermediateValue = memory[287]; /* get 1 */ end
        1106: begin memory[118] = 0; /*set 1 */ end
        1107: begin intermediateValue = memory[292]; /* get 1 */ end
        1108: begin memory[108] = 0; /*set 1 */ end
        1109: begin intermediateValue = memory[293]; /* get 1 */ end
        1110: begin memory[112] = 0; /*set 1 */ end
        1111: begin intermediateValue = memory[294]; /* get 1 */ end
        1112: begin memory[117] = 0; /*set 1 */ end
        1113: begin intermediateValue = memory[289]; /* get 1 */ end
        1114: begin memory[107] = 0; /*set 1 */ end
        1115: begin step =   end.instruction-1; end
        1116: begin intermediateValue = memory[287]; /* get 1 */ end
        1117: begin memory[283] = 0; /*set 1 */ end
        1118: begin memory[114] = 0; /* clear 1 */ end
        1119: begin intermediateValue = memory[283]; /* get 1 */ end
        1120: begin memory[348] = 0; /*set 1 */ end
        1121: begin intermediateValue = memory[113]; /* get 1 */ end
        1122: begin memory[294] = 0; /*set 1 */ end
        1123: begin memory[292] = 0; /*set 1 */ end
        1124: begin memory[293] = 0; /*set 1 */ end
        1125: begin intermediateValue = memory[5]; /* get 2 */ end
        1126: begin memory[344] = 0; /*set 1 */ end
        1127: begin intermediateValue = memory[344]; /* get 1 */ end
        1128: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1129: begin memory[344] = 0; /*set 1 */ end
        1130: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
        1131: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        1132: begin intermediateValue = memory[294]; < memory[166]; ? -1 : memory[294]; == memory[166]; ?  0 : +1; /* compare 2 */ end
        1133: begin if (intermediateValue >  0) step =   end.instruction-1; end
        1134: begin memory[292] = 1; /*set 1 */ end
        1135: begin intermediateValue = memory[166]; /* get 3 */ end
        1136: begin memory[294] = 0; /*set 1 */ end
        1137: begin intermediateValue = memory[25]; /* get 3 */ end
        1138: begin memory[289] = 0; /*set 1 */ end
        1139: begin step =   end.instruction-1; end
        1140: begin intermediateValue = memory[293]; /* get 1 */ end
        1141: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1142: begin memory[293] = 0; /*set 1 */ end
        1143: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
        1144: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        1145: begin step = start.instruction-1; end
        1146: begin intermediateValue = memory[166]; /* get 3 */ end
        1147: begin memory[294] = 0; /*set 1 */ end
        1148: begin intermediateValue = memory[25]; /* get 3 */ end
        1149: begin memory[289] = 0; /*set 1 */ end
        1150: begin intermediateValue = memory[289]; /* get 1 */ end
        1151: begin memory[4] = 0; /*set 1 */ end
        1152: begin intermediateValue = memory[4]; /* get 1 */ end
        1153: begin memory[142] = 0; /*set 1 */ end
        1154: begin intermediateValue = memory[145]; /* get 2 */ end
        1155: begin memory[142] = 0; /*set 1 */ end
        1156: begin intermediateValue = memory[142]; /* get 1 */ end
        1157: begin if (intermediateValue == 0) step =   end.instruction-1; end
        1158: begin intermediateValue = memory[4]; /* get 1 */ end
        1159: begin memory[348] = 0; /*set 1 */ end
        1160: begin intermediateValue = memory[113]; /* get 1 */ end
        1161: begin memory[294] = 0; /*set 1 */ end
        1162: begin memory[292] = 0; /*set 1 */ end
        1163: begin memory[293] = 0; /*set 1 */ end
        1164: begin intermediateValue = memory[5]; /* get 2 */ end
        1165: begin memory[344] = 0; /*set 1 */ end
        1166: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
        1167: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        1168: begin intermediateValue = memory[294]; < memory[166]; ? -1 : memory[294]; == memory[166]; ?  0 : +1; /* compare 2 */ end
        1169: begin if (intermediateValue != 0) step =   end.instruction-1; end
        1170: begin memory[292] = 1; /*set 1 */ end
        1171: begin intermediateValue = memory[166]; /* get 3 */ end
        1172: begin memory[294] = 0; /*set 1 */ end
        1173: begin intermediateValue = memory[25]; /* get 3 */ end
        1174: begin memory[289] = 0; /*set 1 */ end
        1175: begin step =   end.instruction-1; end
        1176: begin intermediateValue = memory[293]; /* get 1 */ end
        1177: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1178: begin memory[293] = 0; /*set 1 */ end
        1179: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
        1180: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        1181: begin step = start.instruction-1; end
        1182: begin intermediateValue = memory[4]; /* get 1 */ end
        1183: begin memory[115] = 0; /*set 1 */ end
        1184: begin intermediateValue = memory[115]; /* get 1 */ end
        1185: begin memory[118] = 0; /*set 1 */ end
        1186: begin intermediateValue = memory[292]; /* get 1 */ end
        1187: begin memory[108] = 0; /*set 1 */ end
        1188: begin intermediateValue = memory[293]; /* get 1 */ end
        1189: begin memory[112] = 0; /*set 1 */ end
        1190: begin intermediateValue = memory[294]; /* get 1 */ end
        1191: begin memory[117] = 0; /*set 1 */ end
        1192: begin intermediateValue = memory[289]; /* get 1 */ end
        1193: begin memory[107] = 0; /*set 1 */ end
        1194: begin step =   end.instruction-1; end
        1195: begin intermediateValue = memory[4]; /* get 1 */ end
        1196: begin memory[283] = 0; /*set 1 */ end
        1197: begin intermediateValue = memory[114]; /* get 1 */ end
        1198: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1199: begin memory[114] = 0; /*set 1 */ end
        1200: begin intermediateValue = memory[114]; /* get 1 */ end
        1201: begin intermediateValue = 9 <  intermediateValue ? -1 : 9 == intermediateValue ?  0 : +1; /* compare 1 */ end
        1202: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        1203: begin step = start.instruction-1; end
        1204: begin $finish("Search did not terminate in a leaf"); end
        1205: begin intermediateValue = memory[108]; /* get 1 */ end
        1206: begin if (intermediateValue == 0) step =   end.instruction-1; end
        1207: begin intermediateValue = memory[118]; /* get 1 */ end
        1208: begin memory[348] = 0; /*set 1 */ end
        1209: begin intermediateValue = memory[111]; /* get 1 */ end
        1210: begin memory[294] = 0; /*set 1 */ end
        1211: begin intermediateValue = memory[110]; /* get 1 */ end
        1212: begin memory[289] = 0; /*set 1 */ end
        1213: begin intermediateValue = memory[112]; /* get 1 */ end
        1214: begin memory[293] = 0; /*set 1 */ end
        1215: begin intermediateValue = memory[294]; /* get 1 */ end
        1216: begin memory[166] = 0; /*set 3 */ end
        1217: begin intermediateValue = memory[289]; /* get 1 */ end
        1218: begin memory[25] = 0; /*set 3 */ end
        1219: begin intermediateValue = memory[293]; < memory[5]; ? -1 : memory[293]; == memory[5]; ?  0 : +1; /* compare 2 */ end
        1220: begin if (intermediateValue <  0) step =   end.instruction-1; end
        1221: begin intermediateValue = memory[5]; /* get 2 */ end
        1222: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1223: begin memory[5] = 0; /*set 2 */ end
        1224: begin memory[140] = 1; /*set 1 */ end
        1225: begin memory[116] = 0; /*set 1 */ end
        1226: begin step =   end.instruction-1; end
        1227: begin intermediateValue = memory[118]; /* get 1 */ end
        1228: begin memory[144] = 0; /*set 1 */ end
        1229: begin intermediateValue = memory[144]; /* get 1 */ end
        1230: begin memory[246] = 0; /*set 1 */ end
        1231: begin intermediateValue = memory[5]; /* get 2 */ end
        1232: begin memory[246] = 0; /*set 1 */ end
        1233: begin intermediateValue = memory[246]; /* get 1 */ end
        1234: begin intermediateValue = 2 <  intermediateValue ? -1 : 2 == intermediateValue ?  0 : +1; /* compare 1 */ end
        1235: begin intermediateValue = intermediateValue >= 0 ? 1 : 0; /* ge */ end
        1236: begin memory[144] = 0; /*set 1 */ end
        1237: begin intermediateValue = memory[144]; /* get 1 */ end
        1238: begin if (intermediateValue >  0) step =   end.instruction-1; end
        1239: begin intermediateValue = memory[118]; /* get 1 */ end
        1240: begin memory[348] = 0; /*set 1 */ end
        1241: begin intermediateValue = memory[111]; /* get 1 */ end
        1242: begin memory[294] = 0; /*set 1 */ end
        1243: begin memory[292] = 0; /*set 1 */ end
        1244: begin memory[293] = 0; /*set 1 */ end
        1245: begin intermediateValue = memory[5]; /* get 2 */ end
        1246: begin memory[344] = 0; /*set 1 */ end
        1247: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
        1248: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        1249: begin intermediateValue = memory[294]; < memory[166]; ? -1 : memory[294]; == memory[166]; ?  0 : +1; /* compare 2 */ end
        1250: begin if (intermediateValue >  0) step =   end.instruction-1; end
        1251: begin memory[292] = 1; /*set 1 */ end
        1252: begin intermediateValue = memory[166]; /* get 3 */ end
        1253: begin memory[294] = 0; /*set 1 */ end
        1254: begin intermediateValue = memory[25]; /* get 3 */ end
        1255: begin memory[289] = 0; /*set 1 */ end
        1256: begin step =   end.instruction-1; end
        1257: begin intermediateValue = memory[293]; /* get 1 */ end
        1258: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1259: begin memory[293] = 0; /*set 1 */ end
        1260: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
        1261: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        1262: begin step = start.instruction-1; end
        1263: begin intermediateValue = memory[118]; /* get 1 */ end
        1264: begin memory[348] = 0; /*set 1 */ end
        1265: begin intermediateValue = memory[111]; /* get 1 */ end
        1266: begin memory[294] = 0; /*set 1 */ end
        1267: begin intermediateValue = memory[110]; /* get 1 */ end
        1268: begin memory[289] = 0; /*set 1 */ end
        1269: begin intermediateValue = memory[293]; /* get 1 */ end
        1270: begin memory[340] = 0; /*set 1 */ end
        1271: begin intermediateValue = memory[5]; /* get 2 */ end
        1272: begin memory[339] = 0; /*set 1 */ end
        1273: begin intermediateValue = memory[339]; /* get 1 */ end
        1274: begin memory[338] = 0; /*set 1 */ end
        1275: begin intermediateValue = memory[338]; /* get 1 */ end
        1276: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1277: begin memory[338] = 0; /*set 1 */ end
        1278: begin intermediateValue = memory[339]; < memory[340]; ? -1 : memory[339]; == memory[340]; ?  0 : +1; /* compare 2 */ end
        1279: begin if (intermediateValue == 0) step =   end.instruction-1; end
        1280: begin intermediateValue = memory[166]; /* get 3 */ end
        1281: begin memory[166] = 0; /*set 3 */ end
        1282: begin intermediateValue = memory[25]; /* get 3 */ end
        1283: begin memory[25] = 0; /*set 3 */ end
        1284: begin intermediateValue = memory[339]; /* get 1 */ end
        1285: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1286: begin memory[339] = 0; /*set 1 */ end
        1287: begin intermediateValue = memory[338]; /* get 1 */ end
        1288: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1289: begin memory[338] = 0; /*set 1 */ end
        1290: begin step = start.instruction-1; end
        1291: begin intermediateValue = memory[294]; /* get 1 */ end
        1292: begin memory[166] = 0; /*set 3 */ end
        1293: begin intermediateValue = memory[289]; /* get 1 */ end
        1294: begin memory[25] = 0; /*set 3 */ end
        1295: begin intermediateValue = memory[5]; /* get 2 */ end
        1296: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1297: begin memory[5] = 0; /*set 2 */ end
        1298: begin memory[140] = 1; /*set 1 */ end
        1299: begin memory[116] = 0; /*set 1 */ end
        1300: begin step =   end.instruction-1; end
        1301: begin memory[140] = 0; /*set 1 */ end
        1302: begin memory[116] = 0; /*set 1 */ end
        1303: begin intermediateValue = memory[285]; /* get 1 */ end
        1304: begin memory[249] = 0; /*set 1 */ end
        1305: begin intermediateValue = memory[145]; /* get 2 */ end
        1306: begin memory[288] = 0; /*set 1 */ end
        1307: begin intermediateValue = memory[288]; /* get 1 */ end
        1308: begin if (intermediateValue >  0) step =   end.instruction-1; end
        1309: begin memory[3] = 0; /* clear 1 */ end
        1310: begin intermediateValue = memory[5]; /* get 2 */ end
        1311: begin memory[3] = 0; /*set 1 */ end
        1312: begin intermediateValue = memory[3]; /* get 1 */ end
        1313: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1314: begin memory[3] = 0; /*set 1 */ end
        1315: begin intermediateValue = memory[3]; /* get 1 */ end
        1316: begin memory[279] = 0; /*set 1 */ end
        1317: begin intermediateValue = memory[279]; /* get 1 */ end
        1318: begin intermediateValue = 1 <  intermediateValue ? -1 : 1 == intermediateValue ?  0 : +1; /* compare 1 */ end
        1319: begin if (intermediateValue >  0) step =   end.instruction-1; end
        1320: begin memory[348] = 0; /*set 1 */ end
        1321: begin memory[293] = 0; /*set 1 */ end
        1322: begin intermediateValue = memory[166]; /* get 3 */ end
        1323: begin memory[294] = 0; /*set 1 */ end
        1324: begin intermediateValue = memory[25]; /* get 3 */ end
        1325: begin memory[289] = 0; /*set 1 */ end
        1326: begin intermediateValue = memory[289]; /* get 1 */ end
        1327: begin memory[276] = 0; /*set 1 */ end
        1328: begin intermediateValue = memory[5]; /* get 2 */ end
        1329: begin memory[293] = 0; /*set 1 */ end
        1330: begin intermediateValue = memory[293]; /* get 1 */ end
        1331: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1332: begin memory[293] = 0; /*set 1 */ end
        1333: begin intermediateValue = memory[166]; /* get 3 */ end
        1334: begin memory[294] = 0; /*set 1 */ end
        1335: begin intermediateValue = memory[25]; /* get 3 */ end
        1336: begin memory[289] = 0; /*set 1 */ end
        1337: begin intermediateValue = memory[289]; /* get 1 */ end
        1338: begin memory[282] = 0; /*set 1 */ end
        1339: begin intermediateValue = memory[287]; /* get 1 */ end
        1340: begin memory[141] = 0; /*set 1 */ end
        1341: begin intermediateValue = memory[25]; /* get 3 */ end
        1342: begin memory[142] = 0; /*set 1 */ end
        1343: begin intermediateValue = memory[145]; /* get 2 */ end
        1344: begin memory[142] = 0; /*set 1 */ end
        1345: begin intermediateValue = memory[142]; /* get 1 */ end
        1346: begin memory[141] = 0; /*set 1 */ end
        1347: begin intermediateValue = memory[141]; /* get 1 */ end
        1348: begin if (intermediateValue == 0) step =   end.instruction-1; end
        1349: begin intermediateValue = memory[276]; /* get 1 */ end
        1350: begin memory[246] = 0; /*set 1 */ end
        1351: begin intermediateValue = memory[5]; /* get 2 */ end
        1352: begin memory[246] = 0; /*set 1 */ end
        1353: begin intermediateValue = memory[246]; /* get 1 */ end
        1354: begin memory[277] = 0; /*set 1 */ end
        1355: begin intermediateValue = memory[282]; /* get 1 */ end
        1356: begin memory[246] = 0; /*set 1 */ end
        1357: begin intermediateValue = memory[5]; /* get 2 */ end
        1358: begin memory[246] = 0; /*set 1 */ end
        1359: begin intermediateValue = memory[246]; /* get 1 */ end
        1360: begin memory[280] = 0; /*set 1 */ end
        1361: begin intermediateValue = memory[277]; /* get 1 */ end
        1362: begin memory[278] = 0; /*set 1 */ end
        1363: begin intermediateValue  = memory[280]; + memory[278];; /* add2 */ end
        1364: begin memory[278] = 0; /*set 1 */ end
        1365: begin intermediateValue = memory[278]; /* get 1 */ end
        1366: begin intermediateValue = 2 <  intermediateValue ? -1 : 2 == intermediateValue ?  0 : +1; /* compare 1 */ end
        1367: begin if (intermediateValue >  0) step =   end.instruction-1; end
        1368: begin intermediateValue = memory[287]; /* get 1 */ end
        1369: begin memory[348] = 0; /*set 1 */ end
        1370: begin memory[5] = 0; /*set 2 */ end
        1371: begin intermediateValue = memory[277]; /* get 1 */ end
        1372: begin intermediateValue = 0 <  intermediateValue ? -1 : 0 == intermediateValue ?  0 : +1; /* compare 1 */ end
        1373: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        1374: begin intermediateValue = memory[276]; /* get 1 */ end
        1375: begin memory[348] = 0; /*set 1 */ end
        1376: begin memory[293] = 0; /* clear 1 */ end
        1377: begin intermediateValue = memory[166]; /* get 3 */ end
        1378: begin memory[294] = 0; /*set 1 */ end
        1379: begin intermediateValue = memory[25]; /* get 3 */ end
        1380: begin memory[289] = 0; /*set 1 */ end
        1381: begin intermediateValue = memory[5]; /* get 2 */ end
        1382: begin memory[347] = 0; /*set 1 */ end
        1383: begin memory[345] = 0; /*set 1 */ end
        1384: begin memory[346] = 1; /*set 1 */ end
        1385: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
        1386: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        1387: begin intermediateValue = memory[166]; /* get 3 */ end
        1388: begin memory[166] = 0; /*set 3 */ end
        1389: begin intermediateValue = memory[25]; /* get 3 */ end
        1390: begin memory[25] = 0; /*set 3 */ end
        1391: begin intermediateValue = memory[345]; /* get 1 */ end
        1392: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1393: begin memory[345] = 0; /*set 1 */ end
        1394: begin intermediateValue = memory[346]; /* get 1 */ end
        1395: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1396: begin memory[346] = 0; /*set 1 */ end
        1397: begin step = start.instruction-1; end
        1398: begin intermediateValue = memory[5]; /* get 2 */ end
        1399: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1400: begin memory[5] = 0; /*set 2 */ end
        1401: begin intermediateValue = memory[287]; /* get 1 */ end
        1402: begin memory[348] = 0; /*set 1 */ end
        1403: begin intermediateValue = memory[5]; /* get 2 */ end
        1404: begin memory[293] = 0; /*set 1 */ end
        1405: begin intermediateValue = memory[294]; /* get 1 */ end
        1406: begin memory[166] = 0; /*set 3 */ end
        1407: begin intermediateValue = memory[289]; /* get 1 */ end
        1408: begin memory[25] = 0; /*set 3 */ end
        1409: begin intermediateValue = memory[5]; /* get 2 */ end
        1410: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1411: begin memory[5] = 0; /*set 2 */ end
        1412: begin intermediateValue = memory[277]; /* get 1 */ end
        1413: begin intermediateValue = 1 <  intermediateValue ? -1 : 1 == intermediateValue ?  0 : +1; /* compare 1 */ end
        1414: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        1415: begin intermediateValue = memory[276]; /* get 1 */ end
        1416: begin memory[348] = 0; /*set 1 */ end
        1417: begin memory[293] = 0; /* clear 1 */ end
        1418: begin intermediateValue = memory[166]; /* get 3 */ end
        1419: begin memory[294] = 0; /*set 1 */ end
        1420: begin intermediateValue = memory[25]; /* get 3 */ end
        1421: begin memory[289] = 0; /*set 1 */ end
        1422: begin intermediateValue = memory[5]; /* get 2 */ end
        1423: begin memory[347] = 0; /*set 1 */ end
        1424: begin memory[345] = 0; /*set 1 */ end
        1425: begin memory[346] = 1; /*set 1 */ end
        1426: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
        1427: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        1428: begin intermediateValue = memory[166]; /* get 3 */ end
        1429: begin memory[166] = 0; /*set 3 */ end
        1430: begin intermediateValue = memory[25]; /* get 3 */ end
        1431: begin memory[25] = 0; /*set 3 */ end
        1432: begin intermediateValue = memory[345]; /* get 1 */ end
        1433: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1434: begin memory[345] = 0; /*set 1 */ end
        1435: begin intermediateValue = memory[346]; /* get 1 */ end
        1436: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1437: begin memory[346] = 0; /*set 1 */ end
        1438: begin step = start.instruction-1; end
        1439: begin intermediateValue = memory[5]; /* get 2 */ end
        1440: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1441: begin memory[5] = 0; /*set 2 */ end
        1442: begin intermediateValue = memory[287]; /* get 1 */ end
        1443: begin memory[348] = 0; /*set 1 */ end
        1444: begin intermediateValue = memory[5]; /* get 2 */ end
        1445: begin memory[293] = 0; /*set 1 */ end
        1446: begin intermediateValue = memory[294]; /* get 1 */ end
        1447: begin memory[166] = 0; /*set 3 */ end
        1448: begin intermediateValue = memory[289]; /* get 1 */ end
        1449: begin memory[25] = 0; /*set 3 */ end
        1450: begin intermediateValue = memory[5]; /* get 2 */ end
        1451: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1452: begin memory[5] = 0; /*set 2 */ end
        1453: begin intermediateValue = memory[280]; /* get 1 */ end
        1454: begin intermediateValue = 0 <  intermediateValue ? -1 : 0 == intermediateValue ?  0 : +1; /* compare 1 */ end
        1455: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        1456: begin intermediateValue = memory[282]; /* get 1 */ end
        1457: begin memory[348] = 0; /*set 1 */ end
        1458: begin memory[293] = 0; /* clear 1 */ end
        1459: begin intermediateValue = memory[166]; /* get 3 */ end
        1460: begin memory[294] = 0; /*set 1 */ end
        1461: begin intermediateValue = memory[25]; /* get 3 */ end
        1462: begin memory[289] = 0; /*set 1 */ end
        1463: begin intermediateValue = memory[5]; /* get 2 */ end
        1464: begin memory[347] = 0; /*set 1 */ end
        1465: begin memory[345] = 0; /*set 1 */ end
        1466: begin memory[346] = 1; /*set 1 */ end
        1467: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
        1468: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        1469: begin intermediateValue = memory[166]; /* get 3 */ end
        1470: begin memory[166] = 0; /*set 3 */ end
        1471: begin intermediateValue = memory[25]; /* get 3 */ end
        1472: begin memory[25] = 0; /*set 3 */ end
        1473: begin intermediateValue = memory[345]; /* get 1 */ end
        1474: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1475: begin memory[345] = 0; /*set 1 */ end
        1476: begin intermediateValue = memory[346]; /* get 1 */ end
        1477: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1478: begin memory[346] = 0; /*set 1 */ end
        1479: begin step = start.instruction-1; end
        1480: begin intermediateValue = memory[5]; /* get 2 */ end
        1481: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1482: begin memory[5] = 0; /*set 2 */ end
        1483: begin intermediateValue = memory[287]; /* get 1 */ end
        1484: begin memory[348] = 0; /*set 1 */ end
        1485: begin intermediateValue = memory[5]; /* get 2 */ end
        1486: begin memory[293] = 0; /*set 1 */ end
        1487: begin intermediateValue = memory[294]; /* get 1 */ end
        1488: begin memory[166] = 0; /*set 3 */ end
        1489: begin intermediateValue = memory[289]; /* get 1 */ end
        1490: begin memory[25] = 0; /*set 3 */ end
        1491: begin intermediateValue = memory[5]; /* get 2 */ end
        1492: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1493: begin memory[5] = 0; /*set 2 */ end
        1494: begin intermediateValue = memory[280]; /* get 1 */ end
        1495: begin intermediateValue = 1 <  intermediateValue ? -1 : 1 == intermediateValue ?  0 : +1; /* compare 1 */ end
        1496: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        1497: begin intermediateValue = memory[282]; /* get 1 */ end
        1498: begin memory[348] = 0; /*set 1 */ end
        1499: begin memory[293] = 0; /* clear 1 */ end
        1500: begin intermediateValue = memory[166]; /* get 3 */ end
        1501: begin memory[294] = 0; /*set 1 */ end
        1502: begin intermediateValue = memory[25]; /* get 3 */ end
        1503: begin memory[289] = 0; /*set 1 */ end
        1504: begin intermediateValue = memory[5]; /* get 2 */ end
        1505: begin memory[347] = 0; /*set 1 */ end
        1506: begin memory[345] = 0; /*set 1 */ end
        1507: begin memory[346] = 1; /*set 1 */ end
        1508: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
        1509: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        1510: begin intermediateValue = memory[166]; /* get 3 */ end
        1511: begin memory[166] = 0; /*set 3 */ end
        1512: begin intermediateValue = memory[25]; /* get 3 */ end
        1513: begin memory[25] = 0; /*set 3 */ end
        1514: begin intermediateValue = memory[345]; /* get 1 */ end
        1515: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1516: begin memory[345] = 0; /*set 1 */ end
        1517: begin intermediateValue = memory[346]; /* get 1 */ end
        1518: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1519: begin memory[346] = 0; /*set 1 */ end
        1520: begin step = start.instruction-1; end
        1521: begin intermediateValue = memory[5]; /* get 2 */ end
        1522: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1523: begin memory[5] = 0; /*set 2 */ end
        1524: begin intermediateValue = memory[287]; /* get 1 */ end
        1525: begin memory[348] = 0; /*set 1 */ end
        1526: begin intermediateValue = memory[5]; /* get 2 */ end
        1527: begin memory[293] = 0; /*set 1 */ end
        1528: begin intermediateValue = memory[294]; /* get 1 */ end
        1529: begin memory[166] = 0; /*set 3 */ end
        1530: begin intermediateValue = memory[289]; /* get 1 */ end
        1531: begin memory[25] = 0; /*set 3 */ end
        1532: begin intermediateValue = memory[5]; /* get 2 */ end
        1533: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1534: begin memory[5] = 0; /*set 2 */ end
        1535: begin intermediateValue = memory[287]; /* get 1 */ end
        1536: begin memory[291] = 0; /*set 1 */ end
        1537: begin memory[145] = 1; /*set 2 */ end
        1538: begin intermediateValue = memory[276]; /* get 1 */ end
        1539: begin memory[120] = -1; /*set 2 */ end
        1540: begin memory[145] = -1; /*set 2 */ end
        1541: begin memory[5] = -1; /*set 2 */ end
        1542: begin memory[166] = -1; /* clear 2 */ end
        1543: begin memory[167] = -1; /* clear 2 */ end
        1544: begin memory[168] = -1; /* clear 2 */ end
        1545: begin memory[169] = -1; /* clear 2 */ end
        1546: begin memory[25] = -1; /* clear 2 */ end
        1547: begin memory[26] = -1; /* clear 2 */ end
        1548: begin memory[27] = -1; /* clear 2 */ end
        1549: begin memory[28] = -1; /* clear 2 */ end
        1550: begin intermediateValue = memory[119]; /* get 1 */ end
        1551: begin memory[120] = 0; /*set 2 */ end
        1552: begin intermediateValue = memory[276]; /* get 1 */ end
        1553: begin memory[119] = 0; /*set 1 */ end
        1554: begin intermediateValue = memory[282]; /* get 1 */ end
        1555: begin memory[120] = -1; /*set 2 */ end
        1556: begin memory[145] = -1; /*set 2 */ end
        1557: begin memory[5] = -1; /*set 2 */ end
        1558: begin memory[166] = -1; /* clear 2 */ end
        1559: begin memory[167] = -1; /* clear 2 */ end
        1560: begin memory[168] = -1; /* clear 2 */ end
        1561: begin memory[169] = -1; /* clear 2 */ end
        1562: begin memory[25] = -1; /* clear 2 */ end
        1563: begin memory[26] = -1; /* clear 2 */ end
        1564: begin memory[27] = -1; /* clear 2 */ end
        1565: begin memory[28] = -1; /* clear 2 */ end
        1566: begin intermediateValue = memory[119]; /* get 1 */ end
        1567: begin memory[120] = 0; /*set 2 */ end
        1568: begin intermediateValue = memory[282]; /* get 1 */ end
        1569: begin memory[119] = 0; /*set 1 */ end
        1570: begin intermediateValue = memory[141]; /* get 1 */ end
        1571: begin if (intermediateValue >  0) step =   end.instruction-1; end
        1572: begin intermediateValue = memory[276]; /* get 1 */ end
        1573: begin memory[3] = 0; /*set 1 */ end
        1574: begin intermediateValue = memory[5]; /* get 2 */ end
        1575: begin memory[3] = 0; /*set 1 */ end
        1576: begin intermediateValue = memory[3]; /* get 1 */ end
        1577: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1578: begin memory[3] = 0; /*set 1 */ end
        1579: begin intermediateValue = memory[3]; /* get 1 */ end
        1580: begin memory[277] = 0; /*set 1 */ end
        1581: begin intermediateValue = memory[282]; /* get 1 */ end
        1582: begin memory[3] = 0; /*set 1 */ end
        1583: begin intermediateValue = memory[5]; /* get 2 */ end
        1584: begin memory[3] = 0; /*set 1 */ end
        1585: begin intermediateValue = memory[3]; /* get 1 */ end
        1586: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1587: begin memory[3] = 0; /*set 1 */ end
        1588: begin intermediateValue = memory[3]; /* get 1 */ end
        1589: begin memory[280] = 0; /*set 1 */ end
        1590: begin intermediateValue = memory[277]; /* get 1 */ end
        1591: begin memory[278] = 0; /*set 1 */ end
        1592: begin intermediateValue  = memory[280]; + memory[278];; /* add2 */ end
        1593: begin memory[278] = 0; /*set 1 */ end
        1594: begin intermediateValue = memory[278]; /* get 1 */ end
        1595: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1596: begin memory[278] = 0; /*set 1 */ end
        1597: begin intermediateValue = memory[278]; /* get 1 */ end
        1598: begin intermediateValue = 3 <  intermediateValue ? -1 : 3 == intermediateValue ?  0 : +1; /* compare 1 */ end
        1599: begin if (intermediateValue >  0) step =   end.instruction-1; end
        1600: begin intermediateValue = memory[287]; /* get 1 */ end
        1601: begin memory[348] = 0; /*set 1 */ end
        1602: begin memory[293] = 0; /*set 1 */ end
        1603: begin intermediateValue = memory[166]; /* get 3 */ end
        1604: begin memory[294] = 0; /*set 1 */ end
        1605: begin intermediateValue = memory[25]; /* get 3 */ end
        1606: begin memory[289] = 0; /*set 1 */ end
        1607: begin intermediateValue = memory[294]; /* get 1 */ end
        1608: begin memory[281] = 0; /*set 1 */ end
        1609: begin memory[5] = 0; /*set 2 */ end
        1610: begin intermediateValue = memory[277]; /* get 1 */ end
        1611: begin intermediateValue = 0 <  intermediateValue ? -1 : 0 == intermediateValue ?  0 : +1; /* compare 1 */ end
        1612: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        1613: begin intermediateValue = memory[276]; /* get 1 */ end
        1614: begin memory[348] = 0; /*set 1 */ end
        1615: begin memory[293] = 0; /* clear 1 */ end
        1616: begin intermediateValue = memory[166]; /* get 3 */ end
        1617: begin memory[294] = 0; /*set 1 */ end
        1618: begin intermediateValue = memory[25]; /* get 3 */ end
        1619: begin memory[289] = 0; /*set 1 */ end
        1620: begin intermediateValue = memory[5]; /* get 2 */ end
        1621: begin memory[347] = 0; /*set 1 */ end
        1622: begin memory[345] = 0; /*set 1 */ end
        1623: begin memory[346] = 1; /*set 1 */ end
        1624: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
        1625: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        1626: begin intermediateValue = memory[166]; /* get 3 */ end
        1627: begin memory[166] = 0; /*set 3 */ end
        1628: begin intermediateValue = memory[25]; /* get 3 */ end
        1629: begin memory[25] = 0; /*set 3 */ end
        1630: begin intermediateValue = memory[345]; /* get 1 */ end
        1631: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1632: begin memory[345] = 0; /*set 1 */ end
        1633: begin intermediateValue = memory[346]; /* get 1 */ end
        1634: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1635: begin memory[346] = 0; /*set 1 */ end
        1636: begin step = start.instruction-1; end
        1637: begin intermediateValue = memory[5]; /* get 2 */ end
        1638: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1639: begin memory[5] = 0; /*set 2 */ end
        1640: begin intermediateValue = memory[287]; /* get 1 */ end
        1641: begin memory[348] = 0; /*set 1 */ end
        1642: begin intermediateValue = memory[5]; /* get 2 */ end
        1643: begin memory[293] = 0; /*set 1 */ end
        1644: begin intermediateValue = memory[294]; /* get 1 */ end
        1645: begin memory[166] = 0; /*set 3 */ end
        1646: begin intermediateValue = memory[289]; /* get 1 */ end
        1647: begin memory[25] = 0; /*set 3 */ end
        1648: begin intermediateValue = memory[5]; /* get 2 */ end
        1649: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1650: begin memory[5] = 0; /*set 2 */ end
        1651: begin intermediateValue = memory[277]; /* get 1 */ end
        1652: begin intermediateValue = 1 <  intermediateValue ? -1 : 1 == intermediateValue ?  0 : +1; /* compare 1 */ end
        1653: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        1654: begin intermediateValue = memory[276]; /* get 1 */ end
        1655: begin memory[348] = 0; /*set 1 */ end
        1656: begin memory[293] = 0; /* clear 1 */ end
        1657: begin intermediateValue = memory[166]; /* get 3 */ end
        1658: begin memory[294] = 0; /*set 1 */ end
        1659: begin intermediateValue = memory[25]; /* get 3 */ end
        1660: begin memory[289] = 0; /*set 1 */ end
        1661: begin intermediateValue = memory[5]; /* get 2 */ end
        1662: begin memory[347] = 0; /*set 1 */ end
        1663: begin memory[345] = 0; /*set 1 */ end
        1664: begin memory[346] = 1; /*set 1 */ end
        1665: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
        1666: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        1667: begin intermediateValue = memory[166]; /* get 3 */ end
        1668: begin memory[166] = 0; /*set 3 */ end
        1669: begin intermediateValue = memory[25]; /* get 3 */ end
        1670: begin memory[25] = 0; /*set 3 */ end
        1671: begin intermediateValue = memory[345]; /* get 1 */ end
        1672: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1673: begin memory[345] = 0; /*set 1 */ end
        1674: begin intermediateValue = memory[346]; /* get 1 */ end
        1675: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1676: begin memory[346] = 0; /*set 1 */ end
        1677: begin step = start.instruction-1; end
        1678: begin intermediateValue = memory[5]; /* get 2 */ end
        1679: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1680: begin memory[5] = 0; /*set 2 */ end
        1681: begin intermediateValue = memory[287]; /* get 1 */ end
        1682: begin memory[348] = 0; /*set 1 */ end
        1683: begin intermediateValue = memory[5]; /* get 2 */ end
        1684: begin memory[293] = 0; /*set 1 */ end
        1685: begin intermediateValue = memory[294]; /* get 1 */ end
        1686: begin memory[166] = 0; /*set 3 */ end
        1687: begin intermediateValue = memory[289]; /* get 1 */ end
        1688: begin memory[25] = 0; /*set 3 */ end
        1689: begin intermediateValue = memory[5]; /* get 2 */ end
        1690: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1691: begin memory[5] = 0; /*set 2 */ end
        1692: begin intermediateValue = memory[277]; /* get 1 */ end
        1693: begin intermediateValue = 2 <  intermediateValue ? -1 : 2 == intermediateValue ?  0 : +1; /* compare 1 */ end
        1694: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        1695: begin intermediateValue = memory[276]; /* get 1 */ end
        1696: begin memory[348] = 0; /*set 1 */ end
        1697: begin memory[293] = 0; /* clear 1 */ end
        1698: begin intermediateValue = memory[166]; /* get 3 */ end
        1699: begin memory[294] = 0; /*set 1 */ end
        1700: begin intermediateValue = memory[25]; /* get 3 */ end
        1701: begin memory[289] = 0; /*set 1 */ end
        1702: begin intermediateValue = memory[5]; /* get 2 */ end
        1703: begin memory[347] = 0; /*set 1 */ end
        1704: begin memory[345] = 0; /*set 1 */ end
        1705: begin memory[346] = 1; /*set 1 */ end
        1706: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
        1707: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        1708: begin intermediateValue = memory[166]; /* get 3 */ end
        1709: begin memory[166] = 0; /*set 3 */ end
        1710: begin intermediateValue = memory[25]; /* get 3 */ end
        1711: begin memory[25] = 0; /*set 3 */ end
        1712: begin intermediateValue = memory[345]; /* get 1 */ end
        1713: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1714: begin memory[345] = 0; /*set 1 */ end
        1715: begin intermediateValue = memory[346]; /* get 1 */ end
        1716: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1717: begin memory[346] = 0; /*set 1 */ end
        1718: begin step = start.instruction-1; end
        1719: begin intermediateValue = memory[5]; /* get 2 */ end
        1720: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1721: begin memory[5] = 0; /*set 2 */ end
        1722: begin intermediateValue = memory[287]; /* get 1 */ end
        1723: begin memory[348] = 0; /*set 1 */ end
        1724: begin intermediateValue = memory[5]; /* get 2 */ end
        1725: begin memory[293] = 0; /*set 1 */ end
        1726: begin intermediateValue = memory[294]; /* get 1 */ end
        1727: begin memory[166] = 0; /*set 3 */ end
        1728: begin intermediateValue = memory[289]; /* get 1 */ end
        1729: begin memory[25] = 0; /*set 3 */ end
        1730: begin intermediateValue = memory[5]; /* get 2 */ end
        1731: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1732: begin memory[5] = 0; /*set 2 */ end
        1733: begin intermediateValue = memory[276]; /* get 1 */ end
        1734: begin memory[348] = 0; /*set 1 */ end
        1735: begin intermediateValue = memory[5]; /* get 2 */ end
        1736: begin memory[293] = 0; /*set 1 */ end
        1737: begin intermediateValue = memory[293]; /* get 1 */ end
        1738: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1739: begin memory[293] = 0; /*set 1 */ end
        1740: begin intermediateValue = memory[166]; /* get 3 */ end
        1741: begin memory[294] = 0; /*set 1 */ end
        1742: begin intermediateValue = memory[25]; /* get 3 */ end
        1743: begin memory[289] = 0; /*set 1 */ end
        1744: begin intermediateValue = memory[287]; /* get 1 */ end
        1745: begin memory[348] = 0; /*set 1 */ end
        1746: begin intermediateValue = memory[281]; /* get 1 */ end
        1747: begin memory[294] = 0; /*set 1 */ end
        1748: begin intermediateValue = memory[5]; /* get 2 */ end
        1749: begin memory[293] = 0; /*set 1 */ end
        1750: begin intermediateValue = memory[294]; /* get 1 */ end
        1751: begin memory[166] = 0; /*set 3 */ end
        1752: begin intermediateValue = memory[289]; /* get 1 */ end
        1753: begin memory[25] = 0; /*set 3 */ end
        1754: begin intermediateValue = memory[5]; /* get 2 */ end
        1755: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1756: begin memory[5] = 0; /*set 2 */ end
        1757: begin intermediateValue = memory[280]; /* get 1 */ end
        1758: begin intermediateValue = 0 <  intermediateValue ? -1 : 0 == intermediateValue ?  0 : +1; /* compare 1 */ end
        1759: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        1760: begin intermediateValue = memory[282]; /* get 1 */ end
        1761: begin memory[348] = 0; /*set 1 */ end
        1762: begin memory[293] = 0; /* clear 1 */ end
        1763: begin intermediateValue = memory[166]; /* get 3 */ end
        1764: begin memory[294] = 0; /*set 1 */ end
        1765: begin intermediateValue = memory[25]; /* get 3 */ end
        1766: begin memory[289] = 0; /*set 1 */ end
        1767: begin intermediateValue = memory[5]; /* get 2 */ end
        1768: begin memory[347] = 0; /*set 1 */ end
        1769: begin memory[345] = 0; /*set 1 */ end
        1770: begin memory[346] = 1; /*set 1 */ end
        1771: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
        1772: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        1773: begin intermediateValue = memory[166]; /* get 3 */ end
        1774: begin memory[166] = 0; /*set 3 */ end
        1775: begin intermediateValue = memory[25]; /* get 3 */ end
        1776: begin memory[25] = 0; /*set 3 */ end
        1777: begin intermediateValue = memory[345]; /* get 1 */ end
        1778: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1779: begin memory[345] = 0; /*set 1 */ end
        1780: begin intermediateValue = memory[346]; /* get 1 */ end
        1781: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1782: begin memory[346] = 0; /*set 1 */ end
        1783: begin step = start.instruction-1; end
        1784: begin intermediateValue = memory[5]; /* get 2 */ end
        1785: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1786: begin memory[5] = 0; /*set 2 */ end
        1787: begin intermediateValue = memory[287]; /* get 1 */ end
        1788: begin memory[348] = 0; /*set 1 */ end
        1789: begin intermediateValue = memory[5]; /* get 2 */ end
        1790: begin memory[293] = 0; /*set 1 */ end
        1791: begin intermediateValue = memory[294]; /* get 1 */ end
        1792: begin memory[166] = 0; /*set 3 */ end
        1793: begin intermediateValue = memory[289]; /* get 1 */ end
        1794: begin memory[25] = 0; /*set 3 */ end
        1795: begin intermediateValue = memory[5]; /* get 2 */ end
        1796: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1797: begin memory[5] = 0; /*set 2 */ end
        1798: begin intermediateValue = memory[280]; /* get 1 */ end
        1799: begin intermediateValue = 1 <  intermediateValue ? -1 : 1 == intermediateValue ?  0 : +1; /* compare 1 */ end
        1800: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        1801: begin intermediateValue = memory[282]; /* get 1 */ end
        1802: begin memory[348] = 0; /*set 1 */ end
        1803: begin memory[293] = 0; /* clear 1 */ end
        1804: begin intermediateValue = memory[166]; /* get 3 */ end
        1805: begin memory[294] = 0; /*set 1 */ end
        1806: begin intermediateValue = memory[25]; /* get 3 */ end
        1807: begin memory[289] = 0; /*set 1 */ end
        1808: begin intermediateValue = memory[5]; /* get 2 */ end
        1809: begin memory[347] = 0; /*set 1 */ end
        1810: begin memory[345] = 0; /*set 1 */ end
        1811: begin memory[346] = 1; /*set 1 */ end
        1812: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
        1813: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        1814: begin intermediateValue = memory[166]; /* get 3 */ end
        1815: begin memory[166] = 0; /*set 3 */ end
        1816: begin intermediateValue = memory[25]; /* get 3 */ end
        1817: begin memory[25] = 0; /*set 3 */ end
        1818: begin intermediateValue = memory[345]; /* get 1 */ end
        1819: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1820: begin memory[345] = 0; /*set 1 */ end
        1821: begin intermediateValue = memory[346]; /* get 1 */ end
        1822: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1823: begin memory[346] = 0; /*set 1 */ end
        1824: begin step = start.instruction-1; end
        1825: begin intermediateValue = memory[5]; /* get 2 */ end
        1826: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1827: begin memory[5] = 0; /*set 2 */ end
        1828: begin intermediateValue = memory[287]; /* get 1 */ end
        1829: begin memory[348] = 0; /*set 1 */ end
        1830: begin intermediateValue = memory[5]; /* get 2 */ end
        1831: begin memory[293] = 0; /*set 1 */ end
        1832: begin intermediateValue = memory[294]; /* get 1 */ end
        1833: begin memory[166] = 0; /*set 3 */ end
        1834: begin intermediateValue = memory[289]; /* get 1 */ end
        1835: begin memory[25] = 0; /*set 3 */ end
        1836: begin intermediateValue = memory[5]; /* get 2 */ end
        1837: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1838: begin memory[5] = 0; /*set 2 */ end
        1839: begin intermediateValue = memory[280]; /* get 1 */ end
        1840: begin intermediateValue = 2 <  intermediateValue ? -1 : 2 == intermediateValue ?  0 : +1; /* compare 1 */ end
        1841: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        1842: begin intermediateValue = memory[282]; /* get 1 */ end
        1843: begin memory[348] = 0; /*set 1 */ end
        1844: begin memory[293] = 0; /* clear 1 */ end
        1845: begin intermediateValue = memory[166]; /* get 3 */ end
        1846: begin memory[294] = 0; /*set 1 */ end
        1847: begin intermediateValue = memory[25]; /* get 3 */ end
        1848: begin memory[289] = 0; /*set 1 */ end
        1849: begin intermediateValue = memory[5]; /* get 2 */ end
        1850: begin memory[347] = 0; /*set 1 */ end
        1851: begin memory[345] = 0; /*set 1 */ end
        1852: begin memory[346] = 1; /*set 1 */ end
        1853: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
        1854: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        1855: begin intermediateValue = memory[166]; /* get 3 */ end
        1856: begin memory[166] = 0; /*set 3 */ end
        1857: begin intermediateValue = memory[25]; /* get 3 */ end
        1858: begin memory[25] = 0; /*set 3 */ end
        1859: begin intermediateValue = memory[345]; /* get 1 */ end
        1860: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1861: begin memory[345] = 0; /*set 1 */ end
        1862: begin intermediateValue = memory[346]; /* get 1 */ end
        1863: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1864: begin memory[346] = 0; /*set 1 */ end
        1865: begin step = start.instruction-1; end
        1866: begin intermediateValue = memory[5]; /* get 2 */ end
        1867: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1868: begin memory[5] = 0; /*set 2 */ end
        1869: begin intermediateValue = memory[287]; /* get 1 */ end
        1870: begin memory[348] = 0; /*set 1 */ end
        1871: begin intermediateValue = memory[5]; /* get 2 */ end
        1872: begin memory[293] = 0; /*set 1 */ end
        1873: begin intermediateValue = memory[294]; /* get 1 */ end
        1874: begin memory[166] = 0; /*set 3 */ end
        1875: begin intermediateValue = memory[289]; /* get 1 */ end
        1876: begin memory[25] = 0; /*set 3 */ end
        1877: begin intermediateValue = memory[5]; /* get 2 */ end
        1878: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1879: begin memory[5] = 0; /*set 2 */ end
        1880: begin intermediateValue = memory[282]; /* get 1 */ end
        1881: begin memory[348] = 0; /*set 1 */ end
        1882: begin intermediateValue = memory[5]; /* get 2 */ end
        1883: begin memory[293] = 0; /*set 1 */ end
        1884: begin intermediateValue = memory[293]; /* get 1 */ end
        1885: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1886: begin memory[293] = 0; /*set 1 */ end
        1887: begin intermediateValue = memory[166]; /* get 3 */ end
        1888: begin memory[294] = 0; /*set 1 */ end
        1889: begin intermediateValue = memory[25]; /* get 3 */ end
        1890: begin memory[289] = 0; /*set 1 */ end
        1891: begin intermediateValue = memory[287]; /* get 1 */ end
        1892: begin memory[348] = 0; /*set 1 */ end
        1893: begin intermediateValue = memory[287]; /* get 1 */ end
        1894: begin memory[294] = 0; /*set 1 */ end
        1895: begin intermediateValue = memory[5]; /* get 2 */ end
        1896: begin memory[293] = 0; /*set 1 */ end
        1897: begin intermediateValue = memory[294]; /* get 1 */ end
        1898: begin memory[166] = 0; /*set 3 */ end
        1899: begin intermediateValue = memory[289]; /* get 1 */ end
        1900: begin memory[25] = 0; /*set 3 */ end
        1901: begin intermediateValue = memory[5]; /* get 2 */ end
        1902: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1903: begin memory[5] = 0; /*set 2 */ end
        1904: begin intermediateValue = memory[276]; /* get 1 */ end
        1905: begin memory[120] = -1; /*set 2 */ end
        1906: begin memory[145] = -1; /*set 2 */ end
        1907: begin memory[5] = -1; /*set 2 */ end
        1908: begin memory[166] = -1; /* clear 2 */ end
        1909: begin memory[167] = -1; /* clear 2 */ end
        1910: begin memory[168] = -1; /* clear 2 */ end
        1911: begin memory[169] = -1; /* clear 2 */ end
        1912: begin memory[25] = -1; /* clear 2 */ end
        1913: begin memory[26] = -1; /* clear 2 */ end
        1914: begin memory[27] = -1; /* clear 2 */ end
        1915: begin memory[28] = -1; /* clear 2 */ end
        1916: begin intermediateValue = memory[119]; /* get 1 */ end
        1917: begin memory[120] = 0; /*set 2 */ end
        1918: begin intermediateValue = memory[276]; /* get 1 */ end
        1919: begin memory[119] = 0; /*set 1 */ end
        1920: begin intermediateValue = memory[282]; /* get 1 */ end
        1921: begin memory[120] = -1; /*set 2 */ end
        1922: begin memory[145] = -1; /*set 2 */ end
        1923: begin memory[5] = -1; /*set 2 */ end
        1924: begin memory[166] = -1; /* clear 2 */ end
        1925: begin memory[167] = -1; /* clear 2 */ end
        1926: begin memory[168] = -1; /* clear 2 */ end
        1927: begin memory[169] = -1; /* clear 2 */ end
        1928: begin memory[25] = -1; /* clear 2 */ end
        1929: begin memory[26] = -1; /* clear 2 */ end
        1930: begin memory[27] = -1; /* clear 2 */ end
        1931: begin memory[28] = -1; /* clear 2 */ end
        1932: begin intermediateValue = memory[119]; /* get 1 */ end
        1933: begin memory[120] = 0; /*set 2 */ end
        1934: begin intermediateValue = memory[282]; /* get 1 */ end
        1935: begin memory[119] = 0; /*set 1 */ end
        1936: begin intermediateValue = memory[287]; /* get 1 */ end
        1937: begin memory[283] = 0; /*set 1 */ end
        1938: begin memory[261] = 0; /* clear 1 */ end
        1939: begin memory[261] = 0; /*set 1 */ end
        1940: begin intermediateValue = memory[283]; /* get 1 */ end
        1941: begin memory[142] = 0; /*set 1 */ end
        1942: begin intermediateValue = memory[145]; /* get 2 */ end
        1943: begin memory[142] = 0; /*set 1 */ end
        1944: begin intermediateValue = memory[142]; /* get 1 */ end
        1945: begin if (intermediateValue >  0) step =   end.instruction-1; end
        1946: begin intermediateValue = memory[283]; /* get 1 */ end
        1947: begin memory[3] = 0; /*set 1 */ end
        1948: begin intermediateValue = memory[5]; /* get 2 */ end
        1949: begin memory[3] = 0; /*set 1 */ end
        1950: begin intermediateValue = memory[3]; /* get 1 */ end
        1951: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1952: begin memory[3] = 0; /*set 1 */ end
        1953: begin intermediateValue = memory[3]; /* get 1 */ end
        1954: begin memory[247] = 0; /*set 1 */ end
        1955: begin intermediateValue = memory[247]; /* get 1 */ end
        1956: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        1957: begin memory[247] = 0; /*set 1 */ end
        1958: begin memory[248] = 0; /*set 1 */ end
        1959: begin intermediateValue = memory[248]; < memory[247]; ? -1 : memory[248]; == memory[247]; ?  0 : +1; /* compare 2 */ end
        1960: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        1961: begin intermediateValue = memory[283]; /* get 1 */ end
        1962: begin memory[256] = 0; /*set 1 */ end
        1963: begin intermediateValue = memory[248]; /* get 1 */ end
        1964: begin memory[251] = 0; /*set 1 */ end
        1965: begin memory[260] = 0; /* clear 1 */ end
        1966: begin intermediateValue = memory[251]; /* get 1 */ end
        1967: begin if (intermediateValue == 0) step =   end.instruction-1; end
        1968: begin intermediateValue = memory[256]; /* get 1 */ end
        1969: begin memory[3] = 0; /*set 1 */ end
        1970: begin intermediateValue = memory[5]; /* get 2 */ end
        1971: begin memory[3] = 0; /*set 1 */ end
        1972: begin intermediateValue = memory[3]; /* get 1 */ end
        1973: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1974: begin memory[3] = 0; /*set 1 */ end
        1975: begin intermediateValue = memory[3]; /* get 1 */ end
        1976: begin memory[250] = 0; /*set 1 */ end
        1977: begin intermediateValue = memory[251]; < memory[250]; ? -1 : memory[251]; == memory[250]; ?  0 : +1; /* compare 2 */ end
        1978: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        1979: begin intermediateValue = memory[256]; /* get 1 */ end
        1980: begin memory[348] = 0; /*set 1 */ end
        1981: begin intermediateValue = memory[251]; /* get 1 */ end
        1982: begin memory[293] = 0; /*set 1 */ end
        1983: begin intermediateValue = memory[293]; /* get 1 */ end
        1984: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        1985: begin memory[293] = 0; /*set 1 */ end
        1986: begin intermediateValue = memory[166]; /* get 3 */ end
        1987: begin memory[294] = 0; /*set 1 */ end
        1988: begin intermediateValue = memory[25]; /* get 3 */ end
        1989: begin memory[289] = 0; /*set 1 */ end
        1990: begin intermediateValue = memory[289]; /* get 1 */ end
        1991: begin memory[252] = 0; /*set 1 */ end
        1992: begin intermediateValue = memory[251]; /* get 1 */ end
        1993: begin memory[293] = 0; /*set 1 */ end
        1994: begin intermediateValue = memory[166]; /* get 3 */ end
        1995: begin memory[294] = 0; /*set 1 */ end
        1996: begin intermediateValue = memory[25]; /* get 3 */ end
        1997: begin memory[289] = 0; /*set 1 */ end
        1998: begin intermediateValue = memory[289]; /* get 1 */ end
        1999: begin memory[257] = 0; /*set 1 */ end
        2000: begin intermediateValue = memory[256]; /* get 1 */ end
        2001: begin memory[141] = 0; /*set 1 */ end
        2002: begin intermediateValue = memory[25]; /* get 3 */ end
        2003: begin memory[142] = 0; /*set 1 */ end
        2004: begin intermediateValue = memory[145]; /* get 2 */ end
        2005: begin memory[142] = 0; /*set 1 */ end
        2006: begin intermediateValue = memory[142]; /* get 1 */ end
        2007: begin memory[141] = 0; /*set 1 */ end
        2008: begin intermediateValue = memory[141]; /* get 1 */ end
        2009: begin if (intermediateValue == 0) step =   end.instruction-1; end
        2010: begin intermediateValue = memory[252]; /* get 1 */ end
        2011: begin memory[246] = 0; /*set 1 */ end
        2012: begin intermediateValue = memory[5]; /* get 2 */ end
        2013: begin memory[246] = 0; /*set 1 */ end
        2014: begin intermediateValue = memory[246]; /* get 1 */ end
        2015: begin memory[253] = 0; /*set 1 */ end
        2016: begin intermediateValue = memory[257]; /* get 1 */ end
        2017: begin memory[246] = 0; /*set 1 */ end
        2018: begin intermediateValue = memory[5]; /* get 2 */ end
        2019: begin memory[246] = 0; /*set 1 */ end
        2020: begin intermediateValue = memory[246]; /* get 1 */ end
        2021: begin memory[255] = 0; /*set 1 */ end
        2022: begin intermediateValue = memory[253]; /* get 1 */ end
        2023: begin memory[254] = 0; /*set 1 */ end
        2024: begin intermediateValue  = memory[255]; + memory[254];; /* add2 */ end
        2025: begin memory[254] = 0; /*set 1 */ end
        2026: begin intermediateValue = memory[254]; /* get 1 */ end
        2027: begin intermediateValue = 2 <  intermediateValue ? -1 : 2 == intermediateValue ?  0 : +1; /* compare 1 */ end
        2028: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        2029: begin intermediateValue = memory[5]; /* get 2 */ end
        2030: begin memory[258] = 0; /*set 1 */ end
        2031: begin intermediateValue = memory[258]; /* get 1 */ end
        2032: begin intermediateValue = 0 <  intermediateValue ? -1 : 0 == intermediateValue ?  0 : +1; /* compare 1 */ end
        2033: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        2034: begin intermediateValue = memory[252]; /* get 1 */ end
        2035: begin memory[348] = 0; /*set 1 */ end
        2036: begin intermediateValue = memory[5]; /* get 2 */ end
        2037: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2038: begin memory[5] = 0; /*set 2 */ end
        2039: begin intermediateValue = memory[5]; /* get 2 */ end
        2040: begin memory[293] = 0; /*set 1 */ end
        2041: begin intermediateValue = memory[166]; /* get 3 */ end
        2042: begin memory[294] = 0; /*set 1 */ end
        2043: begin intermediateValue = memory[25]; /* get 3 */ end
        2044: begin memory[289] = 0; /*set 1 */ end
        2045: begin intermediateValue = memory[257]; /* get 1 */ end
        2046: begin memory[348] = 0; /*set 1 */ end
        2047: begin intermediateValue = memory[5]; /* get 2 */ end
        2048: begin memory[349] = 0; /*set 1 */ end
        2049: begin intermediateValue = memory[349]; /* get 1 */ end
        2050: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        2051: begin intermediateValue = memory[349]; /* get 1 */ end
        2052: begin memory[350] = 0; /*set 1 */ end
        2053: begin intermediateValue = memory[350]; /* get 1 */ end
        2054: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2055: begin memory[350] = 0; /*set 1 */ end
        2056: begin intermediateValue = memory[166]; /* get 3 */ end
        2057: begin memory[166] = 0; /*set 3 */ end
        2058: begin intermediateValue = memory[25]; /* get 3 */ end
        2059: begin memory[25] = 0; /*set 3 */ end
        2060: begin intermediateValue = memory[349]; /* get 1 */ end
        2061: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2062: begin memory[349] = 0; /*set 1 */ end
        2063: begin step = start.instruction-1; end
        2064: begin memory[293] = 0; /*set 1 */ end
        2065: begin intermediateValue = memory[294]; /* get 1 */ end
        2066: begin memory[166] = 0; /*set 3 */ end
        2067: begin intermediateValue = memory[289]; /* get 1 */ end
        2068: begin memory[25] = 0; /*set 3 */ end
        2069: begin intermediateValue = memory[5]; /* get 2 */ end
        2070: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2071: begin memory[5] = 0; /*set 2 */ end
        2072: begin intermediateValue = memory[258]; /* get 1 */ end
        2073: begin intermediateValue = 1 <  intermediateValue ? -1 : 1 == intermediateValue ?  0 : +1; /* compare 1 */ end
        2074: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        2075: begin intermediateValue = memory[252]; /* get 1 */ end
        2076: begin memory[348] = 0; /*set 1 */ end
        2077: begin intermediateValue = memory[5]; /* get 2 */ end
        2078: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2079: begin memory[5] = 0; /*set 2 */ end
        2080: begin intermediateValue = memory[5]; /* get 2 */ end
        2081: begin memory[293] = 0; /*set 1 */ end
        2082: begin intermediateValue = memory[166]; /* get 3 */ end
        2083: begin memory[294] = 0; /*set 1 */ end
        2084: begin intermediateValue = memory[25]; /* get 3 */ end
        2085: begin memory[289] = 0; /*set 1 */ end
        2086: begin intermediateValue = memory[257]; /* get 1 */ end
        2087: begin memory[348] = 0; /*set 1 */ end
        2088: begin intermediateValue = memory[5]; /* get 2 */ end
        2089: begin memory[349] = 0; /*set 1 */ end
        2090: begin intermediateValue = memory[349]; /* get 1 */ end
        2091: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        2092: begin intermediateValue = memory[349]; /* get 1 */ end
        2093: begin memory[350] = 0; /*set 1 */ end
        2094: begin intermediateValue = memory[350]; /* get 1 */ end
        2095: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2096: begin memory[350] = 0; /*set 1 */ end
        2097: begin intermediateValue = memory[166]; /* get 3 */ end
        2098: begin memory[166] = 0; /*set 3 */ end
        2099: begin intermediateValue = memory[25]; /* get 3 */ end
        2100: begin memory[25] = 0; /*set 3 */ end
        2101: begin intermediateValue = memory[349]; /* get 1 */ end
        2102: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2103: begin memory[349] = 0; /*set 1 */ end
        2104: begin step = start.instruction-1; end
        2105: begin memory[293] = 0; /*set 1 */ end
        2106: begin intermediateValue = memory[294]; /* get 1 */ end
        2107: begin memory[166] = 0; /*set 3 */ end
        2108: begin intermediateValue = memory[289]; /* get 1 */ end
        2109: begin memory[25] = 0; /*set 3 */ end
        2110: begin intermediateValue = memory[5]; /* get 2 */ end
        2111: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2112: begin memory[5] = 0; /*set 2 */ end
        2113: begin intermediateValue = memory[141]; /* get 1 */ end
        2114: begin if (intermediateValue >  0) step =   end.instruction-1; end
        2115: begin intermediateValue = memory[252]; /* get 1 */ end
        2116: begin memory[3] = 0; /*set 1 */ end
        2117: begin intermediateValue = memory[5]; /* get 2 */ end
        2118: begin memory[3] = 0; /*set 1 */ end
        2119: begin intermediateValue = memory[3]; /* get 1 */ end
        2120: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2121: begin memory[3] = 0; /*set 1 */ end
        2122: begin intermediateValue = memory[3]; /* get 1 */ end
        2123: begin memory[253] = 0; /*set 1 */ end
        2124: begin intermediateValue = memory[257]; /* get 1 */ end
        2125: begin memory[3] = 0; /*set 1 */ end
        2126: begin intermediateValue = memory[5]; /* get 2 */ end
        2127: begin memory[3] = 0; /*set 1 */ end
        2128: begin intermediateValue = memory[3]; /* get 1 */ end
        2129: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2130: begin memory[3] = 0; /*set 1 */ end
        2131: begin intermediateValue = memory[3]; /* get 1 */ end
        2132: begin memory[255] = 0; /*set 1 */ end
        2133: begin intermediateValue = memory[253]; /* get 1 */ end
        2134: begin memory[254] = 0; /*set 1 */ end
        2135: begin intermediateValue = memory[254]; /* get 1 */ end
        2136: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2137: begin memory[254] = 0; /*set 1 */ end
        2138: begin intermediateValue  = memory[255]; + memory[254];; /* add2 */ end
        2139: begin memory[254] = 0; /*set 1 */ end
        2140: begin intermediateValue = memory[254]; /* get 1 */ end
        2141: begin intermediateValue = 3 <  intermediateValue ? -1 : 3 == intermediateValue ?  0 : +1; /* compare 1 */ end
        2142: begin if (intermediateValue >  0) step =   end.instruction-1; end
        2143: begin intermediateValue = memory[256]; /* get 1 */ end
        2144: begin memory[348] = 0; /*set 1 */ end
        2145: begin intermediateValue = memory[251]; /* get 1 */ end
        2146: begin memory[293] = 0; /*set 1 */ end
        2147: begin intermediateValue = memory[293]; /* get 1 */ end
        2148: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2149: begin memory[293] = 0; /*set 1 */ end
        2150: begin intermediateValue = memory[166]; /* get 3 */ end
        2151: begin memory[294] = 0; /*set 1 */ end
        2152: begin intermediateValue = memory[25]; /* get 3 */ end
        2153: begin memory[289] = 0; /*set 1 */ end
        2154: begin intermediateValue = memory[294]; /* get 1 */ end
        2155: begin memory[259] = 0; /*set 1 */ end
        2156: begin intermediateValue = memory[252]; /* get 1 */ end
        2157: begin memory[348] = 0; /*set 1 */ end
        2158: begin intermediateValue = memory[5]; /* get 2 */ end
        2159: begin memory[293] = 0; /*set 1 */ end
        2160: begin intermediateValue = memory[293]; /* get 1 */ end
        2161: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2162: begin memory[293] = 0; /*set 1 */ end
        2163: begin intermediateValue = memory[166]; /* get 3 */ end
        2164: begin memory[294] = 0; /*set 1 */ end
        2165: begin intermediateValue = memory[25]; /* get 3 */ end
        2166: begin memory[289] = 0; /*set 1 */ end
        2167: begin intermediateValue = memory[257]; /* get 1 */ end
        2168: begin memory[348] = 0; /*set 1 */ end
        2169: begin intermediateValue = memory[259]; /* get 1 */ end
        2170: begin memory[294] = 0; /*set 1 */ end
        2171: begin intermediateValue = memory[5]; /* get 2 */ end
        2172: begin memory[349] = 0; /*set 1 */ end
        2173: begin intermediateValue = memory[349]; /* get 1 */ end
        2174: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        2175: begin intermediateValue = memory[349]; /* get 1 */ end
        2176: begin memory[350] = 0; /*set 1 */ end
        2177: begin intermediateValue = memory[350]; /* get 1 */ end
        2178: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2179: begin memory[350] = 0; /*set 1 */ end
        2180: begin intermediateValue = memory[166]; /* get 3 */ end
        2181: begin memory[166] = 0; /*set 3 */ end
        2182: begin intermediateValue = memory[25]; /* get 3 */ end
        2183: begin memory[25] = 0; /*set 3 */ end
        2184: begin intermediateValue = memory[349]; /* get 1 */ end
        2185: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2186: begin memory[349] = 0; /*set 1 */ end
        2187: begin step = start.instruction-1; end
        2188: begin memory[293] = 0; /*set 1 */ end
        2189: begin intermediateValue = memory[294]; /* get 1 */ end
        2190: begin memory[166] = 0; /*set 3 */ end
        2191: begin intermediateValue = memory[289]; /* get 1 */ end
        2192: begin memory[25] = 0; /*set 3 */ end
        2193: begin intermediateValue = memory[5]; /* get 2 */ end
        2194: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2195: begin memory[5] = 0; /*set 2 */ end
        2196: begin intermediateValue = memory[252]; /* get 1 */ end
        2197: begin memory[348] = 0; /*set 1 */ end
        2198: begin intermediateValue = memory[5]; /* get 2 */ end
        2199: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2200: begin memory[5] = 0; /*set 2 */ end
        2201: begin intermediateValue = memory[5]; /* get 2 */ end
        2202: begin memory[293] = 0; /*set 1 */ end
        2203: begin intermediateValue = memory[166]; /* get 3 */ end
        2204: begin memory[294] = 0; /*set 1 */ end
        2205: begin intermediateValue = memory[25]; /* get 3 */ end
        2206: begin memory[289] = 0; /*set 1 */ end
        2207: begin intermediateValue = memory[252]; /* get 1 */ end
        2208: begin memory[3] = 0; /*set 1 */ end
        2209: begin intermediateValue = memory[5]; /* get 2 */ end
        2210: begin memory[3] = 0; /*set 1 */ end
        2211: begin intermediateValue = memory[3]; /* get 1 */ end
        2212: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2213: begin memory[3] = 0; /*set 1 */ end
        2214: begin intermediateValue = memory[3]; /* get 1 */ end
        2215: begin memory[258] = 0; /*set 1 */ end
        2216: begin intermediateValue = memory[258]; /* get 1 */ end
        2217: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2218: begin memory[258] = 0; /*set 1 */ end
        2219: begin intermediateValue = memory[258]; /* get 1 */ end
        2220: begin intermediateValue = 0 <  intermediateValue ? -1 : 0 == intermediateValue ?  0 : +1; /* compare 1 */ end
        2221: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        2222: begin intermediateValue = memory[252]; /* get 1 */ end
        2223: begin memory[348] = 0; /*set 1 */ end
        2224: begin intermediateValue = memory[5]; /* get 2 */ end
        2225: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2226: begin memory[5] = 0; /*set 2 */ end
        2227: begin intermediateValue = memory[5]; /* get 2 */ end
        2228: begin memory[293] = 0; /*set 1 */ end
        2229: begin intermediateValue = memory[166]; /* get 3 */ end
        2230: begin memory[294] = 0; /*set 1 */ end
        2231: begin intermediateValue = memory[25]; /* get 3 */ end
        2232: begin memory[289] = 0; /*set 1 */ end
        2233: begin intermediateValue = memory[257]; /* get 1 */ end
        2234: begin memory[348] = 0; /*set 1 */ end
        2235: begin intermediateValue = memory[5]; /* get 2 */ end
        2236: begin memory[349] = 0; /*set 1 */ end
        2237: begin intermediateValue = memory[349]; /* get 1 */ end
        2238: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        2239: begin intermediateValue = memory[349]; /* get 1 */ end
        2240: begin memory[350] = 0; /*set 1 */ end
        2241: begin intermediateValue = memory[350]; /* get 1 */ end
        2242: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2243: begin memory[350] = 0; /*set 1 */ end
        2244: begin intermediateValue = memory[166]; /* get 3 */ end
        2245: begin memory[166] = 0; /*set 3 */ end
        2246: begin intermediateValue = memory[25]; /* get 3 */ end
        2247: begin memory[25] = 0; /*set 3 */ end
        2248: begin intermediateValue = memory[349]; /* get 1 */ end
        2249: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2250: begin memory[349] = 0; /*set 1 */ end
        2251: begin step = start.instruction-1; end
        2252: begin memory[293] = 0; /*set 1 */ end
        2253: begin intermediateValue = memory[294]; /* get 1 */ end
        2254: begin memory[166] = 0; /*set 3 */ end
        2255: begin intermediateValue = memory[289]; /* get 1 */ end
        2256: begin memory[25] = 0; /*set 3 */ end
        2257: begin intermediateValue = memory[5]; /* get 2 */ end
        2258: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2259: begin memory[5] = 0; /*set 2 */ end
        2260: begin intermediateValue = memory[258]; /* get 1 */ end
        2261: begin intermediateValue = 1 <  intermediateValue ? -1 : 1 == intermediateValue ?  0 : +1; /* compare 1 */ end
        2262: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        2263: begin intermediateValue = memory[252]; /* get 1 */ end
        2264: begin memory[348] = 0; /*set 1 */ end
        2265: begin intermediateValue = memory[5]; /* get 2 */ end
        2266: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2267: begin memory[5] = 0; /*set 2 */ end
        2268: begin intermediateValue = memory[5]; /* get 2 */ end
        2269: begin memory[293] = 0; /*set 1 */ end
        2270: begin intermediateValue = memory[166]; /* get 3 */ end
        2271: begin memory[294] = 0; /*set 1 */ end
        2272: begin intermediateValue = memory[25]; /* get 3 */ end
        2273: begin memory[289] = 0; /*set 1 */ end
        2274: begin intermediateValue = memory[257]; /* get 1 */ end
        2275: begin memory[348] = 0; /*set 1 */ end
        2276: begin intermediateValue = memory[5]; /* get 2 */ end
        2277: begin memory[349] = 0; /*set 1 */ end
        2278: begin intermediateValue = memory[349]; /* get 1 */ end
        2279: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        2280: begin intermediateValue = memory[349]; /* get 1 */ end
        2281: begin memory[350] = 0; /*set 1 */ end
        2282: begin intermediateValue = memory[350]; /* get 1 */ end
        2283: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2284: begin memory[350] = 0; /*set 1 */ end
        2285: begin intermediateValue = memory[166]; /* get 3 */ end
        2286: begin memory[166] = 0; /*set 3 */ end
        2287: begin intermediateValue = memory[25]; /* get 3 */ end
        2288: begin memory[25] = 0; /*set 3 */ end
        2289: begin intermediateValue = memory[349]; /* get 1 */ end
        2290: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2291: begin memory[349] = 0; /*set 1 */ end
        2292: begin step = start.instruction-1; end
        2293: begin memory[293] = 0; /*set 1 */ end
        2294: begin intermediateValue = memory[294]; /* get 1 */ end
        2295: begin memory[166] = 0; /*set 3 */ end
        2296: begin intermediateValue = memory[289]; /* get 1 */ end
        2297: begin memory[25] = 0; /*set 3 */ end
        2298: begin intermediateValue = memory[5]; /* get 2 */ end
        2299: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2300: begin memory[5] = 0; /*set 2 */ end
        2301: begin intermediateValue = memory[258]; /* get 1 */ end
        2302: begin intermediateValue = 2 <  intermediateValue ? -1 : 2 == intermediateValue ?  0 : +1; /* compare 1 */ end
        2303: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        2304: begin intermediateValue = memory[252]; /* get 1 */ end
        2305: begin memory[348] = 0; /*set 1 */ end
        2306: begin intermediateValue = memory[5]; /* get 2 */ end
        2307: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2308: begin memory[5] = 0; /*set 2 */ end
        2309: begin intermediateValue = memory[5]; /* get 2 */ end
        2310: begin memory[293] = 0; /*set 1 */ end
        2311: begin intermediateValue = memory[166]; /* get 3 */ end
        2312: begin memory[294] = 0; /*set 1 */ end
        2313: begin intermediateValue = memory[25]; /* get 3 */ end
        2314: begin memory[289] = 0; /*set 1 */ end
        2315: begin intermediateValue = memory[257]; /* get 1 */ end
        2316: begin memory[348] = 0; /*set 1 */ end
        2317: begin intermediateValue = memory[5]; /* get 2 */ end
        2318: begin memory[349] = 0; /*set 1 */ end
        2319: begin intermediateValue = memory[349]; /* get 1 */ end
        2320: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        2321: begin intermediateValue = memory[349]; /* get 1 */ end
        2322: begin memory[350] = 0; /*set 1 */ end
        2323: begin intermediateValue = memory[350]; /* get 1 */ end
        2324: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2325: begin memory[350] = 0; /*set 1 */ end
        2326: begin intermediateValue = memory[166]; /* get 3 */ end
        2327: begin memory[166] = 0; /*set 3 */ end
        2328: begin intermediateValue = memory[25]; /* get 3 */ end
        2329: begin memory[25] = 0; /*set 3 */ end
        2330: begin intermediateValue = memory[349]; /* get 1 */ end
        2331: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2332: begin memory[349] = 0; /*set 1 */ end
        2333: begin step = start.instruction-1; end
        2334: begin memory[293] = 0; /*set 1 */ end
        2335: begin intermediateValue = memory[294]; /* get 1 */ end
        2336: begin memory[166] = 0; /*set 3 */ end
        2337: begin intermediateValue = memory[289]; /* get 1 */ end
        2338: begin memory[25] = 0; /*set 3 */ end
        2339: begin intermediateValue = memory[5]; /* get 2 */ end
        2340: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2341: begin memory[5] = 0; /*set 2 */ end
        2342: begin intermediateValue = memory[252]; /* get 1 */ end
        2343: begin memory[120] = -1; /*set 2 */ end
        2344: begin memory[145] = -1; /*set 2 */ end
        2345: begin memory[5] = -1; /*set 2 */ end
        2346: begin memory[166] = -1; /* clear 2 */ end
        2347: begin memory[167] = -1; /* clear 2 */ end
        2348: begin memory[168] = -1; /* clear 2 */ end
        2349: begin memory[169] = -1; /* clear 2 */ end
        2350: begin memory[25] = -1; /* clear 2 */ end
        2351: begin memory[26] = -1; /* clear 2 */ end
        2352: begin memory[27] = -1; /* clear 2 */ end
        2353: begin memory[28] = -1; /* clear 2 */ end
        2354: begin intermediateValue = memory[119]; /* get 1 */ end
        2355: begin memory[120] = 0; /*set 2 */ end
        2356: begin intermediateValue = memory[252]; /* get 1 */ end
        2357: begin memory[119] = 0; /*set 1 */ end
        2358: begin intermediateValue = memory[256]; /* get 1 */ end
        2359: begin memory[348] = 0; /*set 1 */ end
        2360: begin intermediateValue = memory[251]; /* get 1 */ end
        2361: begin memory[293] = 0; /*set 1 */ end
        2362: begin intermediateValue = memory[293]; /* get 1 */ end
        2363: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2364: begin memory[293] = 0; /*set 1 */ end
        2365: begin intermediateValue = memory[5]; /* get 2 */ end
        2366: begin memory[343] = 0; /*set 1 */ end
        2367: begin intermediateValue = memory[293]; /* get 1 */ end
        2368: begin memory[342] = 0; /*set 1 */ end
        2369: begin intermediateValue = memory[342]; /* get 1 */ end
        2370: begin memory[341] = 0; /*set 1 */ end
        2371: begin intermediateValue = memory[341]; /* get 1 */ end
        2372: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2373: begin memory[341] = 0; /*set 1 */ end
        2374: begin intermediateValue = memory[166]; /* get 3 */ end
        2375: begin memory[294] = 0; /*set 1 */ end
        2376: begin intermediateValue = memory[25]; /* get 3 */ end
        2377: begin memory[289] = 0; /*set 1 */ end
        2378: begin intermediateValue = memory[341]; < memory[343]; ? -1 : memory[341]; == memory[343]; ?  0 : +1; /* compare 2 */ end
        2379: begin if (intermediateValue == 0) step =   end.instruction-1; end
        2380: begin intermediateValue = memory[166]; /* get 3 */ end
        2381: begin memory[166] = 0; /*set 3 */ end
        2382: begin intermediateValue = memory[25]; /* get 3 */ end
        2383: begin memory[25] = 0; /*set 3 */ end
        2384: begin intermediateValue = memory[342]; /* get 1 */ end
        2385: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2386: begin memory[342] = 0; /*set 1 */ end
        2387: begin intermediateValue = memory[341]; /* get 1 */ end
        2388: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2389: begin memory[341] = 0; /*set 1 */ end
        2390: begin step = start.instruction-1; end
        2391: begin intermediateValue = memory[5]; /* get 2 */ end
        2392: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2393: begin memory[5] = 0; /*set 2 */ end
        2394: begin memory[260] = 1; /* clear 1 */ end
        2395: begin intermediateValue = memory[260]; /* get 1 */ end
        2396: begin if (intermediateValue == 0) step =   end.instruction-1; end
        2397: begin intermediateValue = memory[248]; /* get 1 */ end
        2398: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2399: begin memory[248] = 0; /*set 1 */ end
        2400: begin intermediateValue = memory[283]; /* get 1 */ end
        2401: begin memory[270] = 0; /*set 1 */ end
        2402: begin intermediateValue = memory[248]; /* get 1 */ end
        2403: begin memory[264] = 0; /*set 1 */ end
        2404: begin memory[275] = 0; /* clear 1 */ end
        2405: begin intermediateValue = memory[5]; /* get 2 */ end
        2406: begin memory[262] = 0; /*set 1 */ end
        2407: begin intermediateValue = memory[262]; /* get 1 */ end
        2408: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2409: begin memory[262] = 0; /*set 1 */ end
        2410: begin intermediateValue = memory[264]; < memory[262]; ? -1 : memory[264]; == memory[262]; ?  0 : +1; /* compare 2 */ end
        2411: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        2412: begin intermediateValue = memory[270]; /* get 1 */ end
        2413: begin memory[348] = 0; /*set 1 */ end
        2414: begin intermediateValue = memory[264]; /* get 1 */ end
        2415: begin memory[293] = 0; /*set 1 */ end
        2416: begin intermediateValue = memory[166]; /* get 3 */ end
        2417: begin memory[294] = 0; /*set 1 */ end
        2418: begin intermediateValue = memory[25]; /* get 3 */ end
        2419: begin memory[289] = 0; /*set 1 */ end
        2420: begin intermediateValue = memory[289]; /* get 1 */ end
        2421: begin memory[266] = 0; /*set 1 */ end
        2422: begin intermediateValue = memory[264]; /* get 1 */ end
        2423: begin memory[293] = 0; /*set 1 */ end
        2424: begin intermediateValue = memory[293]; /* get 1 */ end
        2425: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2426: begin memory[293] = 0; /*set 1 */ end
        2427: begin intermediateValue = memory[166]; /* get 3 */ end
        2428: begin memory[294] = 0; /*set 1 */ end
        2429: begin intermediateValue = memory[25]; /* get 3 */ end
        2430: begin memory[289] = 0; /*set 1 */ end
        2431: begin intermediateValue = memory[289]; /* get 1 */ end
        2432: begin memory[272] = 0; /*set 1 */ end
        2433: begin intermediateValue = memory[270]; /* get 1 */ end
        2434: begin memory[141] = 0; /*set 1 */ end
        2435: begin intermediateValue = memory[25]; /* get 3 */ end
        2436: begin memory[142] = 0; /*set 1 */ end
        2437: begin intermediateValue = memory[145]; /* get 2 */ end
        2438: begin memory[142] = 0; /*set 1 */ end
        2439: begin intermediateValue = memory[142]; /* get 1 */ end
        2440: begin memory[141] = 0; /*set 1 */ end
        2441: begin intermediateValue = memory[141]; /* get 1 */ end
        2442: begin if (intermediateValue == 0) step =   end.instruction-1; end
        2443: begin intermediateValue = memory[266]; /* get 1 */ end
        2444: begin memory[246] = 0; /*set 1 */ end
        2445: begin intermediateValue = memory[5]; /* get 2 */ end
        2446: begin memory[246] = 0; /*set 1 */ end
        2447: begin intermediateValue = memory[246]; /* get 1 */ end
        2448: begin memory[267] = 0; /*set 1 */ end
        2449: begin intermediateValue = memory[272]; /* get 1 */ end
        2450: begin memory[246] = 0; /*set 1 */ end
        2451: begin intermediateValue = memory[5]; /* get 2 */ end
        2452: begin memory[246] = 0; /*set 1 */ end
        2453: begin intermediateValue = memory[246]; /* get 1 */ end
        2454: begin memory[269] = 0; /*set 1 */ end
        2455: begin intermediateValue = memory[267]; /* get 1 */ end
        2456: begin memory[268] = 0; /*set 1 */ end
        2457: begin intermediateValue  = memory[269]; + memory[268];; /* add2 */ end
        2458: begin memory[268] = 0; /*set 1 */ end
        2459: begin intermediateValue = memory[268]; /* get 1 */ end
        2460: begin intermediateValue = 2 <  intermediateValue ? -1 : 2 == intermediateValue ?  0 : +1; /* compare 1 */ end
        2461: begin if (intermediateValue >  0) step =   end.instruction-1; end
        2462: begin intermediateValue = memory[5]; /* get 2 */ end
        2463: begin memory[273] = 0; /*set 1 */ end
        2464: begin intermediateValue = memory[273]; /* get 1 */ end
        2465: begin intermediateValue = 0 <  intermediateValue ? -1 : 0 == intermediateValue ?  0 : +1; /* compare 1 */ end
        2466: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        2467: begin intermediateValue = memory[272]; /* get 1 */ end
        2468: begin memory[348] = 0; /*set 1 */ end
        2469: begin memory[293] = 0; /* clear 1 */ end
        2470: begin intermediateValue = memory[166]; /* get 3 */ end
        2471: begin memory[294] = 0; /*set 1 */ end
        2472: begin intermediateValue = memory[25]; /* get 3 */ end
        2473: begin memory[289] = 0; /*set 1 */ end
        2474: begin intermediateValue = memory[5]; /* get 2 */ end
        2475: begin memory[347] = 0; /*set 1 */ end
        2476: begin memory[345] = 0; /*set 1 */ end
        2477: begin memory[346] = 1; /*set 1 */ end
        2478: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
        2479: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        2480: begin intermediateValue = memory[166]; /* get 3 */ end
        2481: begin memory[166] = 0; /*set 3 */ end
        2482: begin intermediateValue = memory[25]; /* get 3 */ end
        2483: begin memory[25] = 0; /*set 3 */ end
        2484: begin intermediateValue = memory[345]; /* get 1 */ end
        2485: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2486: begin memory[345] = 0; /*set 1 */ end
        2487: begin intermediateValue = memory[346]; /* get 1 */ end
        2488: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2489: begin memory[346] = 0; /*set 1 */ end
        2490: begin step = start.instruction-1; end
        2491: begin intermediateValue = memory[5]; /* get 2 */ end
        2492: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2493: begin memory[5] = 0; /*set 2 */ end
        2494: begin intermediateValue = memory[266]; /* get 1 */ end
        2495: begin memory[348] = 0; /*set 1 */ end
        2496: begin intermediateValue = memory[5]; /* get 2 */ end
        2497: begin memory[293] = 0; /*set 1 */ end
        2498: begin intermediateValue = memory[294]; /* get 1 */ end
        2499: begin memory[166] = 0; /*set 3 */ end
        2500: begin intermediateValue = memory[289]; /* get 1 */ end
        2501: begin memory[25] = 0; /*set 3 */ end
        2502: begin intermediateValue = memory[5]; /* get 2 */ end
        2503: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2504: begin memory[5] = 0; /*set 2 */ end
        2505: begin intermediateValue = memory[273]; /* get 1 */ end
        2506: begin intermediateValue = 1 <  intermediateValue ? -1 : 1 == intermediateValue ?  0 : +1; /* compare 1 */ end
        2507: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        2508: begin intermediateValue = memory[272]; /* get 1 */ end
        2509: begin memory[348] = 0; /*set 1 */ end
        2510: begin memory[293] = 0; /* clear 1 */ end
        2511: begin intermediateValue = memory[166]; /* get 3 */ end
        2512: begin memory[294] = 0; /*set 1 */ end
        2513: begin intermediateValue = memory[25]; /* get 3 */ end
        2514: begin memory[289] = 0; /*set 1 */ end
        2515: begin intermediateValue = memory[5]; /* get 2 */ end
        2516: begin memory[347] = 0; /*set 1 */ end
        2517: begin memory[345] = 0; /*set 1 */ end
        2518: begin memory[346] = 1; /*set 1 */ end
        2519: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
        2520: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        2521: begin intermediateValue = memory[166]; /* get 3 */ end
        2522: begin memory[166] = 0; /*set 3 */ end
        2523: begin intermediateValue = memory[25]; /* get 3 */ end
        2524: begin memory[25] = 0; /*set 3 */ end
        2525: begin intermediateValue = memory[345]; /* get 1 */ end
        2526: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2527: begin memory[345] = 0; /*set 1 */ end
        2528: begin intermediateValue = memory[346]; /* get 1 */ end
        2529: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2530: begin memory[346] = 0; /*set 1 */ end
        2531: begin step = start.instruction-1; end
        2532: begin intermediateValue = memory[5]; /* get 2 */ end
        2533: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2534: begin memory[5] = 0; /*set 2 */ end
        2535: begin intermediateValue = memory[266]; /* get 1 */ end
        2536: begin memory[348] = 0; /*set 1 */ end
        2537: begin intermediateValue = memory[5]; /* get 2 */ end
        2538: begin memory[293] = 0; /*set 1 */ end
        2539: begin intermediateValue = memory[294]; /* get 1 */ end
        2540: begin memory[166] = 0; /*set 3 */ end
        2541: begin intermediateValue = memory[289]; /* get 1 */ end
        2542: begin memory[25] = 0; /*set 3 */ end
        2543: begin intermediateValue = memory[5]; /* get 2 */ end
        2544: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2545: begin memory[5] = 0; /*set 2 */ end
        2546: begin intermediateValue = memory[141]; /* get 1 */ end
        2547: begin if (intermediateValue >  0) step =   end.instruction-1; end
        2548: begin intermediateValue = memory[266]; /* get 1 */ end
        2549: begin memory[3] = 0; /*set 1 */ end
        2550: begin intermediateValue = memory[5]; /* get 2 */ end
        2551: begin memory[3] = 0; /*set 1 */ end
        2552: begin intermediateValue = memory[3]; /* get 1 */ end
        2553: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2554: begin memory[3] = 0; /*set 1 */ end
        2555: begin intermediateValue = memory[3]; /* get 1 */ end
        2556: begin memory[267] = 0; /*set 1 */ end
        2557: begin intermediateValue = memory[272]; /* get 1 */ end
        2558: begin memory[3] = 0; /*set 1 */ end
        2559: begin intermediateValue = memory[5]; /* get 2 */ end
        2560: begin memory[3] = 0; /*set 1 */ end
        2561: begin intermediateValue = memory[3]; /* get 1 */ end
        2562: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2563: begin memory[3] = 0; /*set 1 */ end
        2564: begin intermediateValue = memory[3]; /* get 1 */ end
        2565: begin memory[269] = 0; /*set 1 */ end
        2566: begin intermediateValue = memory[267]; /* get 1 */ end
        2567: begin memory[268] = 0; /*set 1 */ end
        2568: begin intermediateValue = memory[268]; /* get 1 */ end
        2569: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2570: begin memory[268] = 0; /*set 1 */ end
        2571: begin intermediateValue  = memory[269]; + memory[268];; /* add2 */ end
        2572: begin memory[268] = 0; /*set 1 */ end
        2573: begin intermediateValue = memory[268]; /* get 1 */ end
        2574: begin intermediateValue = 3 <  intermediateValue ? -1 : 3 == intermediateValue ?  0 : +1; /* compare 1 */ end
        2575: begin if (intermediateValue >  0) step =   end.instruction-1; end
        2576: begin intermediateValue = memory[266]; /* get 1 */ end
        2577: begin memory[348] = 0; /*set 1 */ end
        2578: begin intermediateValue = memory[5]; /* get 2 */ end
        2579: begin memory[293] = 0; /*set 1 */ end
        2580: begin intermediateValue = memory[293]; /* get 1 */ end
        2581: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2582: begin memory[293] = 0; /*set 1 */ end
        2583: begin intermediateValue = memory[166]; /* get 3 */ end
        2584: begin memory[294] = 0; /*set 1 */ end
        2585: begin intermediateValue = memory[25]; /* get 3 */ end
        2586: begin memory[289] = 0; /*set 1 */ end
        2587: begin intermediateValue = memory[289]; /* get 1 */ end
        2588: begin memory[265] = 0; /*set 1 */ end
        2589: begin intermediateValue = memory[270]; /* get 1 */ end
        2590: begin memory[348] = 0; /*set 1 */ end
        2591: begin intermediateValue = memory[264]; /* get 1 */ end
        2592: begin memory[293] = 0; /*set 1 */ end
        2593: begin intermediateValue = memory[166]; /* get 3 */ end
        2594: begin memory[294] = 0; /*set 1 */ end
        2595: begin intermediateValue = memory[25]; /* get 3 */ end
        2596: begin memory[289] = 0; /*set 1 */ end
        2597: begin intermediateValue = memory[266]; /* get 1 */ end
        2598: begin memory[348] = 0; /*set 1 */ end
        2599: begin intermediateValue = memory[265]; /* get 1 */ end
        2600: begin memory[289] = 0; /*set 1 */ end
        2601: begin intermediateValue = memory[267]; /* get 1 */ end
        2602: begin memory[293] = 0; /*set 1 */ end
        2603: begin intermediateValue = memory[294]; /* get 1 */ end
        2604: begin memory[166] = 0; /*set 3 */ end
        2605: begin intermediateValue = memory[289]; /* get 1 */ end
        2606: begin memory[25] = 0; /*set 3 */ end
        2607: begin intermediateValue = memory[293]; < memory[5]; ? -1 : memory[293]; == memory[5]; ?  0 : +1; /* compare 2 */ end
        2608: begin if (intermediateValue <  0) step =   end.instruction-1; end
        2609: begin intermediateValue = memory[5]; /* get 2 */ end
        2610: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2611: begin memory[5] = 0; /*set 2 */ end
        2612: begin intermediateValue = memory[269]; /* get 1 */ end
        2613: begin memory[273] = 0; /*set 1 */ end
        2614: begin intermediateValue = memory[273]; /* get 1 */ end
        2615: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2616: begin memory[273] = 0; /*set 1 */ end
        2617: begin intermediateValue = memory[273]; /* get 1 */ end
        2618: begin intermediateValue = 0 <  intermediateValue ? -1 : 0 == intermediateValue ?  0 : +1; /* compare 1 */ end
        2619: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        2620: begin intermediateValue = memory[272]; /* get 1 */ end
        2621: begin memory[348] = 0; /*set 1 */ end
        2622: begin memory[293] = 0; /* clear 1 */ end
        2623: begin intermediateValue = memory[166]; /* get 3 */ end
        2624: begin memory[294] = 0; /*set 1 */ end
        2625: begin intermediateValue = memory[25]; /* get 3 */ end
        2626: begin memory[289] = 0; /*set 1 */ end
        2627: begin intermediateValue = memory[5]; /* get 2 */ end
        2628: begin memory[347] = 0; /*set 1 */ end
        2629: begin memory[345] = 0; /*set 1 */ end
        2630: begin memory[346] = 1; /*set 1 */ end
        2631: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
        2632: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        2633: begin intermediateValue = memory[166]; /* get 3 */ end
        2634: begin memory[166] = 0; /*set 3 */ end
        2635: begin intermediateValue = memory[25]; /* get 3 */ end
        2636: begin memory[25] = 0; /*set 3 */ end
        2637: begin intermediateValue = memory[345]; /* get 1 */ end
        2638: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2639: begin memory[345] = 0; /*set 1 */ end
        2640: begin intermediateValue = memory[346]; /* get 1 */ end
        2641: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2642: begin memory[346] = 0; /*set 1 */ end
        2643: begin step = start.instruction-1; end
        2644: begin intermediateValue = memory[5]; /* get 2 */ end
        2645: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2646: begin memory[5] = 0; /*set 2 */ end
        2647: begin intermediateValue = memory[266]; /* get 1 */ end
        2648: begin memory[348] = 0; /*set 1 */ end
        2649: begin intermediateValue = memory[5]; /* get 2 */ end
        2650: begin memory[293] = 0; /*set 1 */ end
        2651: begin intermediateValue = memory[294]; /* get 1 */ end
        2652: begin memory[166] = 0; /*set 3 */ end
        2653: begin intermediateValue = memory[289]; /* get 1 */ end
        2654: begin memory[25] = 0; /*set 3 */ end
        2655: begin intermediateValue = memory[5]; /* get 2 */ end
        2656: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2657: begin memory[5] = 0; /*set 2 */ end
        2658: begin intermediateValue = memory[273]; /* get 1 */ end
        2659: begin intermediateValue = 1 <  intermediateValue ? -1 : 1 == intermediateValue ?  0 : +1; /* compare 1 */ end
        2660: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        2661: begin intermediateValue = memory[272]; /* get 1 */ end
        2662: begin memory[348] = 0; /*set 1 */ end
        2663: begin memory[293] = 0; /* clear 1 */ end
        2664: begin intermediateValue = memory[166]; /* get 3 */ end
        2665: begin memory[294] = 0; /*set 1 */ end
        2666: begin intermediateValue = memory[25]; /* get 3 */ end
        2667: begin memory[289] = 0; /*set 1 */ end
        2668: begin intermediateValue = memory[5]; /* get 2 */ end
        2669: begin memory[347] = 0; /*set 1 */ end
        2670: begin memory[345] = 0; /*set 1 */ end
        2671: begin memory[346] = 1; /*set 1 */ end
        2672: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
        2673: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        2674: begin intermediateValue = memory[166]; /* get 3 */ end
        2675: begin memory[166] = 0; /*set 3 */ end
        2676: begin intermediateValue = memory[25]; /* get 3 */ end
        2677: begin memory[25] = 0; /*set 3 */ end
        2678: begin intermediateValue = memory[345]; /* get 1 */ end
        2679: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2680: begin memory[345] = 0; /*set 1 */ end
        2681: begin intermediateValue = memory[346]; /* get 1 */ end
        2682: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2683: begin memory[346] = 0; /*set 1 */ end
        2684: begin step = start.instruction-1; end
        2685: begin intermediateValue = memory[5]; /* get 2 */ end
        2686: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2687: begin memory[5] = 0; /*set 2 */ end
        2688: begin intermediateValue = memory[266]; /* get 1 */ end
        2689: begin memory[348] = 0; /*set 1 */ end
        2690: begin intermediateValue = memory[5]; /* get 2 */ end
        2691: begin memory[293] = 0; /*set 1 */ end
        2692: begin intermediateValue = memory[294]; /* get 1 */ end
        2693: begin memory[166] = 0; /*set 3 */ end
        2694: begin intermediateValue = memory[289]; /* get 1 */ end
        2695: begin memory[25] = 0; /*set 3 */ end
        2696: begin intermediateValue = memory[5]; /* get 2 */ end
        2697: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2698: begin memory[5] = 0; /*set 2 */ end
        2699: begin intermediateValue = memory[273]; /* get 1 */ end
        2700: begin intermediateValue = 2 <  intermediateValue ? -1 : 2 == intermediateValue ?  0 : +1; /* compare 1 */ end
        2701: begin if (intermediateValue <= 0) step =   end.instruction-1; end
        2702: begin intermediateValue = memory[272]; /* get 1 */ end
        2703: begin memory[348] = 0; /*set 1 */ end
        2704: begin memory[293] = 0; /* clear 1 */ end
        2705: begin intermediateValue = memory[166]; /* get 3 */ end
        2706: begin memory[294] = 0; /*set 1 */ end
        2707: begin intermediateValue = memory[25]; /* get 3 */ end
        2708: begin memory[289] = 0; /*set 1 */ end
        2709: begin intermediateValue = memory[5]; /* get 2 */ end
        2710: begin memory[347] = 0; /*set 1 */ end
        2711: begin memory[345] = 0; /*set 1 */ end
        2712: begin memory[346] = 1; /*set 1 */ end
        2713: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
        2714: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        2715: begin intermediateValue = memory[166]; /* get 3 */ end
        2716: begin memory[166] = 0; /*set 3 */ end
        2717: begin intermediateValue = memory[25]; /* get 3 */ end
        2718: begin memory[25] = 0; /*set 3 */ end
        2719: begin intermediateValue = memory[345]; /* get 1 */ end
        2720: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2721: begin memory[345] = 0; /*set 1 */ end
        2722: begin intermediateValue = memory[346]; /* get 1 */ end
        2723: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2724: begin memory[346] = 0; /*set 1 */ end
        2725: begin step = start.instruction-1; end
        2726: begin intermediateValue = memory[5]; /* get 2 */ end
        2727: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2728: begin memory[5] = 0; /*set 2 */ end
        2729: begin intermediateValue = memory[266]; /* get 1 */ end
        2730: begin memory[348] = 0; /*set 1 */ end
        2731: begin intermediateValue = memory[5]; /* get 2 */ end
        2732: begin memory[293] = 0; /*set 1 */ end
        2733: begin intermediateValue = memory[294]; /* get 1 */ end
        2734: begin memory[166] = 0; /*set 3 */ end
        2735: begin intermediateValue = memory[289]; /* get 1 */ end
        2736: begin memory[25] = 0; /*set 3 */ end
        2737: begin intermediateValue = memory[5]; /* get 2 */ end
        2738: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2739: begin memory[5] = 0; /*set 2 */ end
        2740: begin intermediateValue = memory[272]; /* get 1 */ end
        2741: begin memory[120] = -1; /*set 2 */ end
        2742: begin memory[145] = -1; /*set 2 */ end
        2743: begin memory[5] = -1; /*set 2 */ end
        2744: begin memory[166] = -1; /* clear 2 */ end
        2745: begin memory[167] = -1; /* clear 2 */ end
        2746: begin memory[168] = -1; /* clear 2 */ end
        2747: begin memory[169] = -1; /* clear 2 */ end
        2748: begin memory[25] = -1; /* clear 2 */ end
        2749: begin memory[26] = -1; /* clear 2 */ end
        2750: begin memory[27] = -1; /* clear 2 */ end
        2751: begin memory[28] = -1; /* clear 2 */ end
        2752: begin intermediateValue = memory[119]; /* get 1 */ end
        2753: begin memory[120] = 0; /*set 2 */ end
        2754: begin intermediateValue = memory[272]; /* get 1 */ end
        2755: begin memory[119] = 0; /*set 1 */ end
        2756: begin intermediateValue = memory[270]; /* get 1 */ end
        2757: begin memory[348] = 0; /*set 1 */ end
        2758: begin intermediateValue = memory[264]; /* get 1 */ end
        2759: begin memory[293] = 0; /*set 1 */ end
        2760: begin intermediateValue = memory[293]; /* get 1 */ end
        2761: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2762: begin memory[293] = 0; /*set 1 */ end
        2763: begin intermediateValue = memory[166]; /* get 3 */ end
        2764: begin memory[294] = 0; /*set 1 */ end
        2765: begin intermediateValue = memory[25]; /* get 3 */ end
        2766: begin memory[289] = 0; /*set 1 */ end
        2767: begin intermediateValue = memory[294]; /* get 1 */ end
        2768: begin memory[271] = 0; /*set 1 */ end
        2769: begin intermediateValue = memory[264]; /* get 1 */ end
        2770: begin memory[293] = 0; /*set 1 */ end
        2771: begin intermediateValue = memory[166]; /* get 3 */ end
        2772: begin memory[294] = 0; /*set 1 */ end
        2773: begin intermediateValue = memory[25]; /* get 3 */ end
        2774: begin memory[289] = 0; /*set 1 */ end
        2775: begin intermediateValue = memory[271]; /* get 1 */ end
        2776: begin memory[294] = 0; /*set 1 */ end
        2777: begin intermediateValue = memory[264]; /* get 1 */ end
        2778: begin memory[293] = 0; /*set 1 */ end
        2779: begin intermediateValue = memory[294]; /* get 1 */ end
        2780: begin memory[166] = 0; /*set 3 */ end
        2781: begin intermediateValue = memory[289]; /* get 1 */ end
        2782: begin memory[25] = 0; /*set 3 */ end
        2783: begin intermediateValue = memory[293]; < memory[5]; ? -1 : memory[293]; == memory[5]; ?  0 : +1; /* compare 2 */ end
        2784: begin if (intermediateValue <  0) step =   end.instruction-1; end
        2785: begin intermediateValue = memory[5]; /* get 2 */ end
        2786: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2787: begin memory[5] = 0; /*set 2 */ end
        2788: begin intermediateValue = memory[264]; /* get 1 */ end
        2789: begin memory[293] = 0; /*set 1 */ end
        2790: begin intermediateValue = memory[293]; /* get 1 */ end
        2791: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2792: begin memory[293] = 0; /*set 1 */ end
        2793: begin intermediateValue = memory[5]; /* get 2 */ end
        2794: begin memory[343] = 0; /*set 1 */ end
        2795: begin intermediateValue = memory[293]; /* get 1 */ end
        2796: begin memory[342] = 0; /*set 1 */ end
        2797: begin intermediateValue = memory[342]; /* get 1 */ end
        2798: begin memory[341] = 0; /*set 1 */ end
        2799: begin intermediateValue = memory[341]; /* get 1 */ end
        2800: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2801: begin memory[341] = 0; /*set 1 */ end
        2802: begin intermediateValue = memory[166]; /* get 3 */ end
        2803: begin memory[294] = 0; /*set 1 */ end
        2804: begin intermediateValue = memory[25]; /* get 3 */ end
        2805: begin memory[289] = 0; /*set 1 */ end
        2806: begin intermediateValue = memory[341]; < memory[343]; ? -1 : memory[341]; == memory[343]; ?  0 : +1; /* compare 2 */ end
        2807: begin if (intermediateValue == 0) step =   end.instruction-1; end
        2808: begin intermediateValue = memory[166]; /* get 3 */ end
        2809: begin memory[166] = 0; /*set 3 */ end
        2810: begin intermediateValue = memory[25]; /* get 3 */ end
        2811: begin memory[25] = 0; /*set 3 */ end
        2812: begin intermediateValue = memory[342]; /* get 1 */ end
        2813: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2814: begin memory[342] = 0; /*set 1 */ end
        2815: begin intermediateValue = memory[341]; /* get 1 */ end
        2816: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2817: begin memory[341] = 0; /*set 1 */ end
        2818: begin step = start.instruction-1; end
        2819: begin intermediateValue = memory[5]; /* get 2 */ end
        2820: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2821: begin memory[5] = 0; /*set 2 */ end
        2822: begin memory[275] = 1; /* clear 1 */ end
        2823: begin intermediateValue = memory[248]; /* get 1 */ end
        2824: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2825: begin memory[248] = 0; /*set 1 */ end
        2826: begin step = start.instruction-1; end
        2827: begin intermediateValue = memory[283]; /* get 1 */ end
        2828: begin memory[348] = 0; /*set 1 */ end
        2829: begin intermediateValue = memory[249]; /* get 1 */ end
        2830: begin memory[294] = 0; /*set 1 */ end
        2831: begin memory[292] = 0; /*set 1 */ end
        2832: begin memory[293] = 0; /*set 1 */ end
        2833: begin intermediateValue = memory[5]; /* get 2 */ end
        2834: begin memory[344] = 0; /*set 1 */ end
        2835: begin intermediateValue = memory[344]; /* get 1 */ end
        2836: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2837: begin memory[344] = 0; /*set 1 */ end
        2838: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
        2839: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        2840: begin intermediateValue = memory[294]; < memory[166]; ? -1 : memory[294]; == memory[166]; ?  0 : +1; /* compare 2 */ end
        2841: begin if (intermediateValue >  0) step =   end.instruction-1; end
        2842: begin memory[292] = 1; /*set 1 */ end
        2843: begin intermediateValue = memory[166]; /* get 3 */ end
        2844: begin memory[294] = 0; /*set 1 */ end
        2845: begin intermediateValue = memory[25]; /* get 3 */ end
        2846: begin memory[289] = 0; /*set 1 */ end
        2847: begin step =   end.instruction-1; end
        2848: begin intermediateValue = memory[293]; /* get 1 */ end
        2849: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2850: begin memory[293] = 0; /*set 1 */ end
        2851: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
        2852: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        2853: begin step = start.instruction-1; end
        2854: begin intermediateValue = memory[166]; /* get 3 */ end
        2855: begin memory[294] = 0; /*set 1 */ end
        2856: begin intermediateValue = memory[25]; /* get 3 */ end
        2857: begin memory[289] = 0; /*set 1 */ end
        2858: begin intermediateValue = memory[289]; /* get 1 */ end
        2859: begin memory[283] = 0; /*set 1 */ end
        2860: begin intermediateValue = memory[261]; /* get 1 */ end
        2861: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2862: begin memory[261] = 0; /*set 1 */ end
        2863: begin intermediateValue = memory[261]; /* get 1 */ end
        2864: begin intermediateValue = 9 <  intermediateValue ? -1 : 9 == intermediateValue ?  0 : +1; /* compare 1 */ end
        2865: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        2866: begin step = start.instruction-1; end
        2867: begin $finish("Fallen off the end of the tree"); end
        2868: begin step =   end.instruction-1; end
        2869: begin intermediateValue = memory[4]; /* get 1 */ end
        2870: begin memory[144] = 0; /*set 1 */ end
        2871: begin intermediateValue = memory[144]; /* get 1 */ end
        2872: begin memory[3] = 0; /*set 1 */ end
        2873: begin intermediateValue = memory[5]; /* get 2 */ end
        2874: begin memory[3] = 0; /*set 1 */ end
        2875: begin intermediateValue = memory[3]; /* get 1 */ end
        2876: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2877: begin memory[3] = 0; /*set 1 */ end
        2878: begin intermediateValue = memory[3]; /* get 1 */ end
        2879: begin intermediateValue = 3 <  intermediateValue ? -1 : 3 == intermediateValue ?  0 : +1; /* compare 1 */ end
        2880: begin intermediateValue = intermediateValue >= 0 ? 1 : 0; /* ge */ end
        2881: begin memory[144] = 0; /*set 1 */ end
        2882: begin intermediateValue = memory[144]; /* get 1 */ end
        2883: begin if (intermediateValue == 0) step =   end.instruction-1; end
        2884: begin intermediateValue = memory[4]; /* get 1 */ end
        2885: begin memory[297] = 0; /*set 1 */ end
        2886: begin intermediateValue = memory[283]; /* get 1 */ end
        2887: begin memory[298] = 0; /*set 1 */ end
        2888: begin intermediateValue = memory[293]; /* get 1 */ end
        2889: begin memory[295] = 0; /*set 1 */ end
        2890: begin intermediateValue = memory[119]; /* get 1 */ end
        2891: begin memory[296] = 0; /*set 1 */ end
        2892: begin intermediateValue = memory[296]; /* get 1 */ end
        2893: begin if (intermediateValue >  0) step =   end.instruction-1; end
        2894: begin $finish("No more memory available"); end
        2895: begin intermediateValue = memory[120]; /* get 2 */ end
        2896: begin memory[119] = 0; /*set 1 */ end
        2897: begin memory[120] = 0; /*set 2 */ end
        2898: begin memory[145] = 0; /*set 2 */ end
        2899: begin memory[5] = 0; /*set 2 */ end
        2900: begin memory[166] = 0; /* clear 2 */ end
        2901: begin memory[167] = 0; /* clear 2 */ end
        2902: begin memory[168] = 0; /* clear 2 */ end
        2903: begin memory[169] = 0; /* clear 2 */ end
        2904: begin memory[25] = 0; /* clear 2 */ end
        2905: begin memory[26] = 0; /* clear 2 */ end
        2906: begin memory[27] = 0; /* clear 2 */ end
        2907: begin memory[28] = 0; /* clear 2 */ end
        2908: begin intermediateValue = memory[296]; /* get 1 */ end
        2909: begin memory[290] = 0; /*set 1 */ end
        2910: begin memory[145] = 0; /*set 2 */ end
        2911: begin intermediateValue = memory[297]; /* get 1 */ end
        2912: begin memory[348] = 0; /*set 1 */ end
        2913: begin memory[293] = 0; /* clear 1 */ end
        2914: begin intermediateValue = memory[166]; /* get 3 */ end
        2915: begin memory[294] = 0; /*set 1 */ end
        2916: begin intermediateValue = memory[25]; /* get 3 */ end
        2917: begin memory[289] = 0; /*set 1 */ end
        2918: begin intermediateValue = memory[5]; /* get 2 */ end
        2919: begin memory[347] = 0; /*set 1 */ end
        2920: begin memory[345] = 0; /*set 1 */ end
        2921: begin memory[346] = 1; /*set 1 */ end
        2922: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
        2923: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        2924: begin intermediateValue = memory[166]; /* get 3 */ end
        2925: begin memory[166] = 0; /*set 3 */ end
        2926: begin intermediateValue = memory[25]; /* get 3 */ end
        2927: begin memory[25] = 0; /*set 3 */ end
        2928: begin intermediateValue = memory[345]; /* get 1 */ end
        2929: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2930: begin memory[345] = 0; /*set 1 */ end
        2931: begin intermediateValue = memory[346]; /* get 1 */ end
        2932: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2933: begin memory[346] = 0; /*set 1 */ end
        2934: begin step = start.instruction-1; end
        2935: begin intermediateValue = memory[5]; /* get 2 */ end
        2936: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2937: begin memory[5] = 0; /*set 2 */ end
        2938: begin intermediateValue = memory[296]; /* get 1 */ end
        2939: begin memory[348] = 0; /*set 1 */ end
        2940: begin intermediateValue = memory[5]; /* get 2 */ end
        2941: begin memory[293] = 0; /*set 1 */ end
        2942: begin intermediateValue = memory[294]; /* get 1 */ end
        2943: begin memory[166] = 0; /*set 3 */ end
        2944: begin intermediateValue = memory[289]; /* get 1 */ end
        2945: begin memory[25] = 0; /*set 3 */ end
        2946: begin intermediateValue = memory[5]; /* get 2 */ end
        2947: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2948: begin memory[5] = 0; /*set 2 */ end
        2949: begin intermediateValue = memory[297]; /* get 1 */ end
        2950: begin memory[348] = 0; /*set 1 */ end
        2951: begin memory[293] = 0; /* clear 1 */ end
        2952: begin intermediateValue = memory[166]; /* get 3 */ end
        2953: begin memory[294] = 0; /*set 1 */ end
        2954: begin intermediateValue = memory[25]; /* get 3 */ end
        2955: begin memory[289] = 0; /*set 1 */ end
        2956: begin intermediateValue = memory[5]; /* get 2 */ end
        2957: begin memory[347] = 0; /*set 1 */ end
        2958: begin memory[345] = 0; /*set 1 */ end
        2959: begin memory[346] = 1; /*set 1 */ end
        2960: begin intermediateValue = memory[346]; < memory[347]; ? -1 : memory[346]; == memory[347]; ?  0 : +1; /* compare 2 */ end
        2961: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        2962: begin intermediateValue = memory[166]; /* get 3 */ end
        2963: begin memory[166] = 0; /*set 3 */ end
        2964: begin intermediateValue = memory[25]; /* get 3 */ end
        2965: begin memory[25] = 0; /*set 3 */ end
        2966: begin intermediateValue = memory[345]; /* get 1 */ end
        2967: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2968: begin memory[345] = 0; /*set 1 */ end
        2969: begin intermediateValue = memory[346]; /* get 1 */ end
        2970: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2971: begin memory[346] = 0; /*set 1 */ end
        2972: begin step = start.instruction-1; end
        2973: begin intermediateValue = memory[5]; /* get 2 */ end
        2974: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        2975: begin memory[5] = 0; /*set 2 */ end
        2976: begin intermediateValue = memory[294]; /* get 1 */ end
        2977: begin memory[299] = 0; /*set 1 */ end
        2978: begin intermediateValue = memory[296]; /* get 1 */ end
        2979: begin memory[348] = 0; /*set 1 */ end
        2980: begin intermediateValue = memory[287]; /* get 1 */ end
        2981: begin memory[294] = 0; /*set 1 */ end
        2982: begin intermediateValue = memory[5]; /* get 2 */ end
        2983: begin memory[293] = 0; /*set 1 */ end
        2984: begin intermediateValue = memory[294]; /* get 1 */ end
        2985: begin memory[166] = 0; /*set 3 */ end
        2986: begin intermediateValue = memory[289]; /* get 1 */ end
        2987: begin memory[25] = 0; /*set 3 */ end
        2988: begin intermediateValue = memory[5]; /* get 2 */ end
        2989: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        2990: begin memory[5] = 0; /*set 2 */ end
        2991: begin intermediateValue = memory[298]; /* get 1 */ end
        2992: begin memory[348] = 0; /*set 1 */ end
        2993: begin intermediateValue = memory[299]; /* get 1 */ end
        2994: begin memory[294] = 0; /*set 1 */ end
        2995: begin intermediateValue = memory[296]; /* get 1 */ end
        2996: begin memory[289] = 0; /*set 1 */ end
        2997: begin intermediateValue = memory[295]; /* get 1 */ end
        2998: begin memory[293] = 0; /*set 1 */ end
        2999: begin intermediateValue = memory[293]; /* get 1 */ end
        3000: begin memory[340] = 0; /*set 1 */ end
        3001: begin intermediateValue = memory[5]; /* get 2 */ end
        3002: begin memory[339] = 0; /*set 1 */ end
        3003: begin intermediateValue = memory[339]; /* get 1 */ end
        3004: begin memory[338] = 0; /*set 1 */ end
        3005: begin intermediateValue = memory[338]; /* get 1 */ end
        3006: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        3007: begin memory[338] = 0; /*set 1 */ end
        3008: begin intermediateValue = memory[339]; < memory[340]; ? -1 : memory[339]; == memory[340]; ?  0 : +1; /* compare 2 */ end
        3009: begin if (intermediateValue == 0) step =   end.instruction-1; end
        3010: begin intermediateValue = memory[166]; /* get 3 */ end
        3011: begin memory[166] = 0; /*set 3 */ end
        3012: begin intermediateValue = memory[25]; /* get 3 */ end
        3013: begin memory[25] = 0; /*set 3 */ end
        3014: begin intermediateValue = memory[339]; /* get 1 */ end
        3015: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        3016: begin memory[339] = 0; /*set 1 */ end
        3017: begin intermediateValue = memory[338]; /* get 1 */ end
        3018: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        3019: begin memory[338] = 0; /*set 1 */ end
        3020: begin step = start.instruction-1; end
        3021: begin intermediateValue = memory[294]; /* get 1 */ end
        3022: begin memory[166] = 0; /*set 3 */ end
        3023: begin intermediateValue = memory[289]; /* get 1 */ end
        3024: begin memory[25] = 0; /*set 3 */ end
        3025: begin intermediateValue = memory[5]; /* get 2 */ end
        3026: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        3027: begin memory[5] = 0; /*set 2 */ end
        3028: begin intermediateValue = memory[283]; /* get 1 */ end
        3029: begin memory[348] = 0; /*set 1 */ end
        3030: begin intermediateValue = memory[285]; /* get 1 */ end
        3031: begin memory[294] = 0; /*set 1 */ end
        3032: begin memory[292] = 0; /*set 1 */ end
        3033: begin memory[293] = 0; /*set 1 */ end
        3034: begin intermediateValue = memory[5]; /* get 2 */ end
        3035: begin memory[344] = 0; /*set 1 */ end
        3036: begin intermediateValue = memory[344]; /* get 1 */ end
        3037: begin intermediateValue = -1 + intermediateValue;  /* add 1 */ end
        3038: begin memory[344] = 0; /*set 1 */ end
        3039: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
        3040: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        3041: begin intermediateValue = memory[294]; < memory[166]; ? -1 : memory[294]; == memory[166]; ?  0 : +1; /* compare 2 */ end
        3042: begin if (intermediateValue >  0) step =   end.instruction-1; end
        3043: begin memory[292] = 1; /*set 1 */ end
        3044: begin intermediateValue = memory[166]; /* get 3 */ end
        3045: begin memory[294] = 0; /*set 1 */ end
        3046: begin intermediateValue = memory[25]; /* get 3 */ end
        3047: begin memory[289] = 0; /*set 1 */ end
        3048: begin step =   end.instruction-1; end
        3049: begin intermediateValue = memory[293]; /* get 1 */ end
        3050: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        3051: begin memory[293] = 0; /*set 1 */ end
        3052: begin intermediateValue = memory[293]; < memory[344]; ? -1 : memory[293]; == memory[344]; ?  0 : +1; /* compare 2 */ end
        3053: begin if (intermediateValue >= 0) step =   end.instruction-1; end
        3054: begin step = start.instruction-1; end
        3055: begin intermediateValue = memory[166]; /* get 3 */ end
        3056: begin memory[294] = 0; /*set 1 */ end
        3057: begin intermediateValue = memory[25]; /* get 3 */ end
        3058: begin memory[289] = 0; /*set 1 */ end
        3059: begin intermediateValue = memory[289]; /* get 1 */ end
        3060: begin memory[283] = 0; /*set 1 */ end
        3061: begin intermediateValue = memory[144]; /* get 1 */ end
        3062: begin if (intermediateValue >  0) step =   end.instruction-1; end
        3063: begin intermediateValue = memory[4]; /* get 1 */ end
        3064: begin memory[283] = 0; /*set 1 */ end
        3065: begin intermediateValue = memory[286]; /* get 1 */ end
        3066: begin intermediateValue = 1 + intermediateValue;  /* add 1 */ end
        3067: begin memory[286] = 0; /*set 1 */ end
        3068: begin intermediateValue = memory[286]; /* get 1 */ end
        3069: begin intermediateValue = 9 <  intermediateValue ? -1 : 9 == intermediateValue ?  0 : +1; /* compare 1 */ end
        3070: begin if (intermediateValue >  0) step =   end.instruction-1; end
        3071: begin step = start.instruction-1; end
        3072: begin $finish("Fallen off the end of the tree"); end

        endcase
    end // Execute
  end // Always
endmodule
