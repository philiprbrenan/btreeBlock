//-----------------------------------------------------------------------------
// Generic cpu
// Philip R Brenan at appaapps dot com, Appa Apps Ltd Inc., 2025-01-07
//------------------------------------------------------------------------------
`timescale 10ps/1ps
(* keep_hierarchy = "yes" *)
module find(reset, stop, clock, Key, Data, data, found);                    // Database on a chip
  input                      reset;                                             // Restart the program run sequence when this goes high
  input                      clock;                                             // Program counter clock
  input [16-1:0]  Key;                                             // Input key
  input [16-1:0] Data;                                             // Input data
  output                      stop;                                             // Program has stopped when this goes high
  output[16-1:0] data;                                             // Output data
  output                     found;                                             // Whether the key was found on put, find delete

  integer step;
  integer steps;
  integer stopped;
  integer intermediateValue;
  reg [16-1:0] memory [23531-1: 0];


  assign stop  = stopped > 0 ? 1 : 0;
  assign found = memory[11408];
  assign data  = memory[11407];

  always @ (posedge clock) begin                                                // Execute next step in program
    if (reset) begin                                                            // Reset
      step     <= 0;
      steps    <= 0;
      stopped  <= 0;
      begin
        integer i;
        for (i = 0; i < 23531; i = i + 1) begin
          memory[i] <= 0;
        end
      end
      memory[   3] <=   15; /* branchSize */
      memory[   4] <=    2; /* child */
      memory[   5] <=   16; /* current_size[0] */
      memory[   6] <=   16; /* current_size[1] */
      memory[   7] <=   16; /* current_size[2] */
      memory[   8] <=   16; /* current_size[3] */
      memory[   9] <=   16; /* current_size[4] */
      memory[  10] <=   16; /* current_size[5] */
      memory[  11] <=   16; /* current_size[6] */
      memory[  12] <=   16; /* current_size[7] */
      memory[  13] <=   16; /* current_size[8] */
      memory[  14] <=   16; /* current_size[9] */
      memory[  15] <=   16; /* current_size[10] */
      memory[  16] <=   16; /* current_size[11] */
      memory[  17] <=   16; /* current_size[12] */
      memory[  18] <=   16; /* current_size[13] */
      memory[  19] <=   16; /* current_size[14] */
      memory[  20] <=   16; /* current_size[15] */
      memory[  21] <=   16; /* current_size[16] */
      memory[  22] <=   -1; /* current_size[17] */
      memory[ 605] <=    1; /* data[0,0] */
      memory[ 606] <=    3; /* data[0,1] */
      memory[ 607] <=    4; /* data[0,2] */
      memory[ 608] <=    5; /* data[0,3] */
      memory[ 609] <=    6; /* data[0,4] */
      memory[ 610] <=    7; /* data[0,5] */
      memory[ 611] <=    8; /* data[0,6] */
      memory[ 612] <=    9; /* data[0,7] */
      memory[ 613] <=   10; /* data[0,8] */
      memory[ 614] <=   11; /* data[0,9] */
      memory[ 615] <=   12; /* data[0,10] */
      memory[ 616] <=   13; /* data[0,11] */
      memory[ 617] <=   14; /* data[0,12] */
      memory[ 618] <=   15; /* data[0,13] */
      memory[ 619] <=   16; /* data[0,14] */
      memory[ 620] <=    2; /* data[0,15] */
      memory[ 621] <=    2; /* data[0,16] */
      memory[ 623] <=  256; /* data[1,0] */
      memory[ 624] <=  255; /* data[1,1] */
      memory[ 625] <=  254; /* data[1,2] */
      memory[ 626] <=  253; /* data[1,3] */
      memory[ 627] <=  252; /* data[1,4] */
      memory[ 628] <=  251; /* data[1,5] */
      memory[ 629] <=  250; /* data[1,6] */
      memory[ 630] <=  249; /* data[1,7] */
      memory[ 631] <=  248; /* data[1,8] */
      memory[ 632] <=  247; /* data[1,9] */
      memory[ 633] <=  246; /* data[1,10] */
      memory[ 634] <=  245; /* data[1,11] */
      memory[ 635] <=  244; /* data[1,12] */
      memory[ 636] <=  243; /* data[1,13] */
      memory[ 637] <=  242; /* data[1,14] */
      memory[ 638] <=  241; /* data[1,15] */
      memory[ 641] <=   16; /* data[2,0] */
      memory[ 642] <=   15; /* data[2,1] */
      memory[ 643] <=   14; /* data[2,2] */
      memory[ 644] <=   13; /* data[2,3] */
      memory[ 645] <=   12; /* data[2,4] */
      memory[ 646] <=   11; /* data[2,5] */
      memory[ 647] <=   10; /* data[2,6] */
      memory[ 648] <=    9; /* data[2,7] */
      memory[ 649] <=    8; /* data[2,8] */
      memory[ 650] <=    7; /* data[2,9] */
      memory[ 651] <=    6; /* data[2,10] */
      memory[ 652] <=    5; /* data[2,11] */
      memory[ 653] <=    4; /* data[2,12] */
      memory[ 654] <=    3; /* data[2,13] */
      memory[ 655] <=    2; /* data[2,14] */
      memory[ 656] <=    1; /* data[2,15] */
      memory[ 659] <=  240; /* data[3,0] */
      memory[ 660] <=  239; /* data[3,1] */
      memory[ 661] <=  238; /* data[3,2] */
      memory[ 662] <=  237; /* data[3,3] */
      memory[ 663] <=  236; /* data[3,4] */
      memory[ 664] <=  235; /* data[3,5] */
      memory[ 665] <=  234; /* data[3,6] */
      memory[ 666] <=  233; /* data[3,7] */
      memory[ 667] <=  232; /* data[3,8] */
      memory[ 668] <=  231; /* data[3,9] */
      memory[ 669] <=  230; /* data[3,10] */
      memory[ 670] <=  229; /* data[3,11] */
      memory[ 671] <=  228; /* data[3,12] */
      memory[ 672] <=  227; /* data[3,13] */
      memory[ 673] <=  226; /* data[3,14] */
      memory[ 674] <=  225; /* data[3,15] */
      memory[ 677] <=  224; /* data[4,0] */
      memory[ 678] <=  223; /* data[4,1] */
      memory[ 679] <=  222; /* data[4,2] */
      memory[ 680] <=  221; /* data[4,3] */
      memory[ 681] <=  220; /* data[4,4] */
      memory[ 682] <=  219; /* data[4,5] */
      memory[ 683] <=  218; /* data[4,6] */
      memory[ 684] <=  217; /* data[4,7] */
      memory[ 685] <=  216; /* data[4,8] */
      memory[ 686] <=  215; /* data[4,9] */
      memory[ 687] <=  214; /* data[4,10] */
      memory[ 688] <=  213; /* data[4,11] */
      memory[ 689] <=  212; /* data[4,12] */
      memory[ 690] <=  211; /* data[4,13] */
      memory[ 691] <=  210; /* data[4,14] */
      memory[ 692] <=  209; /* data[4,15] */
      memory[ 695] <=  208; /* data[5,0] */
      memory[ 696] <=  207; /* data[5,1] */
      memory[ 697] <=  206; /* data[5,2] */
      memory[ 698] <=  205; /* data[5,3] */
      memory[ 699] <=  204; /* data[5,4] */
      memory[ 700] <=  203; /* data[5,5] */
      memory[ 701] <=  202; /* data[5,6] */
      memory[ 702] <=  201; /* data[5,7] */
      memory[ 703] <=  200; /* data[5,8] */
      memory[ 704] <=  199; /* data[5,9] */
      memory[ 705] <=  198; /* data[5,10] */
      memory[ 706] <=  197; /* data[5,11] */
      memory[ 707] <=  196; /* data[5,12] */
      memory[ 708] <=  195; /* data[5,13] */
      memory[ 709] <=  194; /* data[5,14] */
      memory[ 710] <=  193; /* data[5,15] */
      memory[ 713] <=  192; /* data[6,0] */
      memory[ 714] <=  191; /* data[6,1] */
      memory[ 715] <=  190; /* data[6,2] */
      memory[ 716] <=  189; /* data[6,3] */
      memory[ 717] <=  188; /* data[6,4] */
      memory[ 718] <=  187; /* data[6,5] */
      memory[ 719] <=  186; /* data[6,6] */
      memory[ 720] <=  185; /* data[6,7] */
      memory[ 721] <=  184; /* data[6,8] */
      memory[ 722] <=  183; /* data[6,9] */
      memory[ 723] <=  182; /* data[6,10] */
      memory[ 724] <=  181; /* data[6,11] */
      memory[ 725] <=  180; /* data[6,12] */
      memory[ 726] <=  179; /* data[6,13] */
      memory[ 727] <=  178; /* data[6,14] */
      memory[ 728] <=  177; /* data[6,15] */
      memory[ 731] <=  176; /* data[7,0] */
      memory[ 732] <=  175; /* data[7,1] */
      memory[ 733] <=  174; /* data[7,2] */
      memory[ 734] <=  173; /* data[7,3] */
      memory[ 735] <=  172; /* data[7,4] */
      memory[ 736] <=  171; /* data[7,5] */
      memory[ 737] <=  170; /* data[7,6] */
      memory[ 738] <=  169; /* data[7,7] */
      memory[ 739] <=  168; /* data[7,8] */
      memory[ 740] <=  167; /* data[7,9] */
      memory[ 741] <=  166; /* data[7,10] */
      memory[ 742] <=  165; /* data[7,11] */
      memory[ 743] <=  164; /* data[7,12] */
      memory[ 744] <=  163; /* data[7,13] */
      memory[ 745] <=  162; /* data[7,14] */
      memory[ 746] <=  161; /* data[7,15] */
      memory[ 749] <=  160; /* data[8,0] */
      memory[ 750] <=  159; /* data[8,1] */
      memory[ 751] <=  158; /* data[8,2] */
      memory[ 752] <=  157; /* data[8,3] */
      memory[ 753] <=  156; /* data[8,4] */
      memory[ 754] <=  155; /* data[8,5] */
      memory[ 755] <=  154; /* data[8,6] */
      memory[ 756] <=  153; /* data[8,7] */
      memory[ 757] <=  152; /* data[8,8] */
      memory[ 758] <=  151; /* data[8,9] */
      memory[ 759] <=  150; /* data[8,10] */
      memory[ 760] <=  149; /* data[8,11] */
      memory[ 761] <=  148; /* data[8,12] */
      memory[ 762] <=  147; /* data[8,13] */
      memory[ 763] <=  146; /* data[8,14] */
      memory[ 764] <=  145; /* data[8,15] */
      memory[ 767] <=  144; /* data[9,0] */
      memory[ 768] <=  143; /* data[9,1] */
      memory[ 769] <=  142; /* data[9,2] */
      memory[ 770] <=  141; /* data[9,3] */
      memory[ 771] <=  140; /* data[9,4] */
      memory[ 772] <=  139; /* data[9,5] */
      memory[ 773] <=  138; /* data[9,6] */
      memory[ 774] <=  137; /* data[9,7] */
      memory[ 775] <=  136; /* data[9,8] */
      memory[ 776] <=  135; /* data[9,9] */
      memory[ 777] <=  134; /* data[9,10] */
      memory[ 778] <=  133; /* data[9,11] */
      memory[ 779] <=  132; /* data[9,12] */
      memory[ 780] <=  131; /* data[9,13] */
      memory[ 781] <=  130; /* data[9,14] */
      memory[ 782] <=  129; /* data[9,15] */
      memory[ 785] <=  128; /* data[10,0] */
      memory[ 786] <=  127; /* data[10,1] */
      memory[ 787] <=  126; /* data[10,2] */
      memory[ 788] <=  125; /* data[10,3] */
      memory[ 789] <=  124; /* data[10,4] */
      memory[ 790] <=  123; /* data[10,5] */
      memory[ 791] <=  122; /* data[10,6] */
      memory[ 792] <=  121; /* data[10,7] */
      memory[ 793] <=  120; /* data[10,8] */
      memory[ 794] <=  119; /* data[10,9] */
      memory[ 795] <=  118; /* data[10,10] */
      memory[ 796] <=  117; /* data[10,11] */
      memory[ 797] <=  116; /* data[10,12] */
      memory[ 798] <=  115; /* data[10,13] */
      memory[ 799] <=  114; /* data[10,14] */
      memory[ 800] <=  113; /* data[10,15] */
      memory[ 803] <=  112; /* data[11,0] */
      memory[ 804] <=  111; /* data[11,1] */
      memory[ 805] <=  110; /* data[11,2] */
      memory[ 806] <=  109; /* data[11,3] */
      memory[ 807] <=  108; /* data[11,4] */
      memory[ 808] <=  107; /* data[11,5] */
      memory[ 809] <=  106; /* data[11,6] */
      memory[ 810] <=  105; /* data[11,7] */
      memory[ 811] <=  104; /* data[11,8] */
      memory[ 812] <=  103; /* data[11,9] */
      memory[ 813] <=  102; /* data[11,10] */
      memory[ 814] <=  101; /* data[11,11] */
      memory[ 815] <=  100; /* data[11,12] */
      memory[ 816] <=   99; /* data[11,13] */
      memory[ 817] <=   98; /* data[11,14] */
      memory[ 818] <=   97; /* data[11,15] */
      memory[ 821] <=   96; /* data[12,0] */
      memory[ 822] <=   95; /* data[12,1] */
      memory[ 823] <=   94; /* data[12,2] */
      memory[ 824] <=   93; /* data[12,3] */
      memory[ 825] <=   92; /* data[12,4] */
      memory[ 826] <=   91; /* data[12,5] */
      memory[ 827] <=   90; /* data[12,6] */
      memory[ 828] <=   89; /* data[12,7] */
      memory[ 829] <=   88; /* data[12,8] */
      memory[ 830] <=   87; /* data[12,9] */
      memory[ 831] <=   86; /* data[12,10] */
      memory[ 832] <=   85; /* data[12,11] */
      memory[ 833] <=   84; /* data[12,12] */
      memory[ 834] <=   83; /* data[12,13] */
      memory[ 835] <=   82; /* data[12,14] */
      memory[ 836] <=   81; /* data[12,15] */
      memory[ 839] <=   80; /* data[13,0] */
      memory[ 840] <=   79; /* data[13,1] */
      memory[ 841] <=   78; /* data[13,2] */
      memory[ 842] <=   77; /* data[13,3] */
      memory[ 843] <=   76; /* data[13,4] */
      memory[ 844] <=   75; /* data[13,5] */
      memory[ 845] <=   74; /* data[13,6] */
      memory[ 846] <=   73; /* data[13,7] */
      memory[ 847] <=   72; /* data[13,8] */
      memory[ 848] <=   71; /* data[13,9] */
      memory[ 849] <=   70; /* data[13,10] */
      memory[ 850] <=   69; /* data[13,11] */
      memory[ 851] <=   68; /* data[13,12] */
      memory[ 852] <=   67; /* data[13,13] */
      memory[ 853] <=   66; /* data[13,14] */
      memory[ 854] <=   65; /* data[13,15] */
      memory[ 857] <=   64; /* data[14,0] */
      memory[ 858] <=   63; /* data[14,1] */
      memory[ 859] <=   62; /* data[14,2] */
      memory[ 860] <=   61; /* data[14,3] */
      memory[ 861] <=   60; /* data[14,4] */
      memory[ 862] <=   59; /* data[14,5] */
      memory[ 863] <=   58; /* data[14,6] */
      memory[ 864] <=   57; /* data[14,7] */
      memory[ 865] <=   56; /* data[14,8] */
      memory[ 866] <=   55; /* data[14,9] */
      memory[ 867] <=   54; /* data[14,10] */
      memory[ 868] <=   53; /* data[14,11] */
      memory[ 869] <=   52; /* data[14,12] */
      memory[ 870] <=   51; /* data[14,13] */
      memory[ 871] <=   50; /* data[14,14] */
      memory[ 872] <=   49; /* data[14,15] */
      memory[ 875] <=   48; /* data[15,0] */
      memory[ 876] <=   47; /* data[15,1] */
      memory[ 877] <=   46; /* data[15,2] */
      memory[ 878] <=   45; /* data[15,3] */
      memory[ 879] <=   44; /* data[15,4] */
      memory[ 880] <=   43; /* data[15,5] */
      memory[ 881] <=   42; /* data[15,6] */
      memory[ 882] <=   41; /* data[15,7] */
      memory[ 883] <=   40; /* data[15,8] */
      memory[ 884] <=   39; /* data[15,9] */
      memory[ 885] <=   38; /* data[15,10] */
      memory[ 886] <=   37; /* data[15,11] */
      memory[ 887] <=   36; /* data[15,12] */
      memory[ 888] <=   35; /* data[15,13] */
      memory[ 889] <=   34; /* data[15,14] */
      memory[ 890] <=   33; /* data[15,15] */
      memory[ 893] <=   32; /* data[16,0] */
      memory[ 894] <=   31; /* data[16,1] */
      memory[ 895] <=   30; /* data[16,2] */
      memory[ 896] <=   29; /* data[16,3] */
      memory[ 897] <=   28; /* data[16,4] */
      memory[ 898] <=   27; /* data[16,5] */
      memory[ 899] <=   26; /* data[16,6] */
      memory[ 900] <=   25; /* data[16,7] */
      memory[ 901] <=   24; /* data[16,8] */
      memory[ 902] <=   23; /* data[16,9] */
      memory[ 903] <=   22; /* data[16,10] */
      memory[ 904] <=   21; /* data[16,11] */
      memory[ 905] <=   20; /* data[16,12] */
      memory[ 906] <=   19; /* data[16,13] */
      memory[ 907] <=   18; /* data[16,14] */
      memory[ 908] <=   17; /* data[16,15] */
      memory[ 911] <=   -1; /* data[17,0] */
      memory[ 912] <=   -1; /* data[17,1] */
      memory[ 913] <=   -1; /* data[17,2] */
      memory[ 914] <=   -1; /* data[17,3] */
      memory[ 915] <=   -1; /* data[17,4] */
      memory[ 916] <=   -1; /* data[17,5] */
      memory[ 917] <=   -1; /* data[17,6] */
      memory[ 918] <=   -1; /* data[17,7] */
      memory[ 919] <=   -1; /* data[17,8] */
      memory[ 920] <=   -1; /* data[17,9] */
      memory[ 921] <=   -1; /* data[17,10] */
      memory[ 922] <=   -1; /* data[17,11] */
      memory[ 923] <=   -1; /* data[17,12] */
      memory[ 924] <=   -1; /* data[17,13] */
      memory[ 925] <=   -1; /* data[17,14] */
      memory[ 926] <=   -1; /* data[17,15] */
      memory[ 927] <=   -1; /* data[17,16] */
      memory[ 928] <=   -1; /* data[17,17] */
      memory[11407] <=    2; /* f_data */
      memory[11410] <=    1; /* findAndInsert_Data */
      memory[11411] <=  256; /* findAndInsert_Key */
      memory[11412] <=   15; /* f_index */
      memory[11413] <=  256; /* find_Key */
      memory[11415] <=    2; /* find_result_leaf */
      memory[11417] <=  256; /* f_key */
      memory[11418] <=    2; /* f_leaf */
      memory[11419] <=   17; /* freeChainHead */
      memory[11437] <=   18; /* free[17] */
      memory[11438] <=   19; /* free[18] */
      memory[11439] <=   20; /* free[19] */
      memory[11440] <=   21; /* free[20] */
      memory[11441] <=   22; /* free[21] */
      memory[11442] <=   23; /* free[22] */
      memory[11443] <=   24; /* free[23] */
      memory[11444] <=   25; /* free[24] */
      memory[11445] <=   26; /* free[25] */
      memory[11446] <=   27; /* free[26] */
      memory[11447] <=   28; /* free[27] */
      memory[11448] <=   29; /* free[28] */
      memory[11449] <=   30; /* free[29] */
      memory[11450] <=   31; /* free[30] */
      memory[11451] <=   32; /* free[31] */
      memory[11452] <=   33; /* free[32] */
      memory[11453] <=   34; /* free[33] */
      memory[11454] <=   35; /* free[34] */
      memory[11455] <=   36; /* free[35] */
      memory[11456] <=   37; /* free[36] */
      memory[11457] <=   38; /* free[37] */
      memory[11458] <=   39; /* free[38] */
      memory[11459] <=   40; /* free[39] */
      memory[11460] <=   41; /* free[40] */
      memory[11461] <=   42; /* free[41] */
      memory[11462] <=   43; /* free[42] */
      memory[11463] <=   44; /* free[43] */
      memory[11464] <=   45; /* free[44] */
      memory[11465] <=   46; /* free[45] */
      memory[11466] <=   47; /* free[46] */
      memory[11467] <=   48; /* free[47] */
      memory[11468] <=   49; /* free[48] */
      memory[11469] <=   50; /* free[49] */
      memory[11470] <=   51; /* free[50] */
      memory[11471] <=   52; /* free[51] */
      memory[11472] <=   53; /* free[52] */
      memory[11473] <=   54; /* free[53] */
      memory[11474] <=   55; /* free[54] */
      memory[11475] <=   56; /* free[55] */
      memory[11476] <=   57; /* free[56] */
      memory[11477] <=   58; /* free[57] */
      memory[11478] <=   59; /* free[58] */
      memory[11479] <=   60; /* free[59] */
      memory[11480] <=   61; /* free[60] */
      memory[11481] <=   62; /* free[61] */
      memory[11482] <=   63; /* free[62] */
      memory[11483] <=   64; /* free[63] */
      memory[11484] <=   65; /* free[64] */
      memory[11485] <=   66; /* free[65] */
      memory[11486] <=   67; /* free[66] */
      memory[11487] <=   68; /* free[67] */
      memory[11488] <=   69; /* free[68] */
      memory[11489] <=   70; /* free[69] */
      memory[11490] <=   71; /* free[70] */
      memory[11491] <=   72; /* free[71] */
      memory[11492] <=   73; /* free[72] */
      memory[11493] <=   74; /* free[73] */
      memory[11494] <=   75; /* free[74] */
      memory[11495] <=   76; /* free[75] */
      memory[11496] <=   77; /* free[76] */
      memory[11497] <=   78; /* free[77] */
      memory[11498] <=   79; /* free[78] */
      memory[11499] <=   80; /* free[79] */
      memory[11500] <=   81; /* free[80] */
      memory[11501] <=   82; /* free[81] */
      memory[11502] <=   83; /* free[82] */
      memory[11503] <=   84; /* free[83] */
      memory[11504] <=   85; /* free[84] */
      memory[11505] <=   86; /* free[85] */
      memory[11506] <=   87; /* free[86] */
      memory[11507] <=   88; /* free[87] */
      memory[11508] <=   89; /* free[88] */
      memory[11509] <=   90; /* free[89] */
      memory[11510] <=   91; /* free[90] */
      memory[11511] <=   92; /* free[91] */
      memory[11512] <=   93; /* free[92] */
      memory[11513] <=   94; /* free[93] */
      memory[11514] <=   95; /* free[94] */
      memory[11515] <=   96; /* free[95] */
      memory[11516] <=   97; /* free[96] */
      memory[11517] <=   98; /* free[97] */
      memory[11518] <=   99; /* free[98] */
      memory[11519] <=  100; /* free[99] */
      memory[11520] <=  101; /* free[100] */
      memory[11521] <=  102; /* free[101] */
      memory[11522] <=  103; /* free[102] */
      memory[11523] <=  104; /* free[103] */
      memory[11524] <=  105; /* free[104] */
      memory[11525] <=  106; /* free[105] */
      memory[11526] <=  107; /* free[106] */
      memory[11527] <=  108; /* free[107] */
      memory[11528] <=  109; /* free[108] */
      memory[11529] <=  110; /* free[109] */
      memory[11530] <=  111; /* free[110] */
      memory[11531] <=  112; /* free[111] */
      memory[11532] <=  113; /* free[112] */
      memory[11533] <=  114; /* free[113] */
      memory[11534] <=  115; /* free[114] */
      memory[11535] <=  116; /* free[115] */
      memory[11536] <=  117; /* free[116] */
      memory[11537] <=  118; /* free[117] */
      memory[11538] <=  119; /* free[118] */
      memory[11539] <=  120; /* free[119] */
      memory[11540] <=  121; /* free[120] */
      memory[11541] <=  122; /* free[121] */
      memory[11542] <=  123; /* free[122] */
      memory[11543] <=  124; /* free[123] */
      memory[11544] <=  125; /* free[124] */
      memory[11545] <=  126; /* free[125] */
      memory[11546] <=  127; /* free[126] */
      memory[11547] <=  128; /* free[127] */
      memory[11548] <=  129; /* free[128] */
      memory[11549] <=  130; /* free[129] */
      memory[11550] <=  131; /* free[130] */
      memory[11551] <=  132; /* free[131] */
      memory[11552] <=  133; /* free[132] */
      memory[11553] <=  134; /* free[133] */
      memory[11554] <=  135; /* free[134] */
      memory[11555] <=  136; /* free[135] */
      memory[11556] <=  137; /* free[136] */
      memory[11557] <=  138; /* free[137] */
      memory[11558] <=  139; /* free[138] */
      memory[11559] <=  140; /* free[139] */
      memory[11560] <=  141; /* free[140] */
      memory[11561] <=  142; /* free[141] */
      memory[11562] <=  143; /* free[142] */
      memory[11563] <=  144; /* free[143] */
      memory[11564] <=  145; /* free[144] */
      memory[11565] <=  146; /* free[145] */
      memory[11566] <=  147; /* free[146] */
      memory[11567] <=  148; /* free[147] */
      memory[11568] <=  149; /* free[148] */
      memory[11569] <=  150; /* free[149] */
      memory[11570] <=  151; /* free[150] */
      memory[11571] <=  152; /* free[151] */
      memory[11572] <=  153; /* free[152] */
      memory[11573] <=  154; /* free[153] */
      memory[11574] <=  155; /* free[154] */
      memory[11575] <=  156; /* free[155] */
      memory[11576] <=  157; /* free[156] */
      memory[11577] <=  158; /* free[157] */
      memory[11578] <=  159; /* free[158] */
      memory[11579] <=  160; /* free[159] */
      memory[11580] <=  161; /* free[160] */
      memory[11581] <=  162; /* free[161] */
      memory[11582] <=  163; /* free[162] */
      memory[11583] <=  164; /* free[163] */
      memory[11584] <=  165; /* free[164] */
      memory[11585] <=  166; /* free[165] */
      memory[11586] <=  167; /* free[166] */
      memory[11587] <=  168; /* free[167] */
      memory[11588] <=  169; /* free[168] */
      memory[11589] <=  170; /* free[169] */
      memory[11590] <=  171; /* free[170] */
      memory[11591] <=  172; /* free[171] */
      memory[11592] <=  173; /* free[172] */
      memory[11593] <=  174; /* free[173] */
      memory[11594] <=  175; /* free[174] */
      memory[11595] <=  176; /* free[175] */
      memory[11596] <=  177; /* free[176] */
      memory[11597] <=  178; /* free[177] */
      memory[11598] <=  179; /* free[178] */
      memory[11599] <=  180; /* free[179] */
      memory[11600] <=  181; /* free[180] */
      memory[11601] <=  182; /* free[181] */
      memory[11602] <=  183; /* free[182] */
      memory[11603] <=  184; /* free[183] */
      memory[11604] <=  185; /* free[184] */
      memory[11605] <=  186; /* free[185] */
      memory[11606] <=  187; /* free[186] */
      memory[11607] <=  188; /* free[187] */
      memory[11608] <=  189; /* free[188] */
      memory[11609] <=  190; /* free[189] */
      memory[11610] <=  191; /* free[190] */
      memory[11611] <=  192; /* free[191] */
      memory[11612] <=  193; /* free[192] */
      memory[11613] <=  194; /* free[193] */
      memory[11614] <=  195; /* free[194] */
      memory[11615] <=  196; /* free[195] */
      memory[11616] <=  197; /* free[196] */
      memory[11617] <=  198; /* free[197] */
      memory[11618] <=  199; /* free[198] */
      memory[11619] <=  200; /* free[199] */
      memory[11620] <=  201; /* free[200] */
      memory[11621] <=  202; /* free[201] */
      memory[11622] <=  203; /* free[202] */
      memory[11623] <=  204; /* free[203] */
      memory[11624] <=  205; /* free[204] */
      memory[11625] <=  206; /* free[205] */
      memory[11626] <=  207; /* free[206] */
      memory[11627] <=  208; /* free[207] */
      memory[11628] <=  209; /* free[208] */
      memory[11629] <=  210; /* free[209] */
      memory[11630] <=  211; /* free[210] */
      memory[11631] <=  212; /* free[211] */
      memory[11632] <=  213; /* free[212] */
      memory[11633] <=  214; /* free[213] */
      memory[11634] <=  215; /* free[214] */
      memory[11635] <=  216; /* free[215] */
      memory[11636] <=  217; /* free[216] */
      memory[11637] <=  218; /* free[217] */
      memory[11638] <=  219; /* free[218] */
      memory[11639] <=  220; /* free[219] */
      memory[11640] <=  221; /* free[220] */
      memory[11641] <=  222; /* free[221] */
      memory[11642] <=  223; /* free[222] */
      memory[11643] <=  224; /* free[223] */
      memory[11644] <=  225; /* free[224] */
      memory[11645] <=  226; /* free[225] */
      memory[11646] <=  227; /* free[226] */
      memory[11647] <=  228; /* free[227] */
      memory[11648] <=  229; /* free[228] */
      memory[11649] <=  230; /* free[229] */
      memory[11650] <=  231; /* free[230] */
      memory[11651] <=  232; /* free[231] */
      memory[11652] <=  233; /* free[232] */
      memory[11653] <=  234; /* free[233] */
      memory[11654] <=  235; /* free[234] */
      memory[11655] <=  236; /* free[235] */
      memory[11656] <=  237; /* free[236] */
      memory[11657] <=  238; /* free[237] */
      memory[11658] <=  239; /* free[238] */
      memory[11659] <=  240; /* free[239] */
      memory[11660] <=  241; /* free[240] */
      memory[11661] <=  242; /* free[241] */
      memory[11662] <=  243; /* free[242] */
      memory[11663] <=  244; /* free[243] */
      memory[11664] <=  245; /* free[244] */
      memory[11665] <=  246; /* free[245] */
      memory[11666] <=  247; /* free[246] */
      memory[11667] <=  248; /* free[247] */
      memory[11668] <=  249; /* free[248] */
      memory[11669] <=  250; /* free[249] */
      memory[11670] <=  251; /* free[250] */
      memory[11671] <=  252; /* free[251] */
      memory[11672] <=  253; /* free[252] */
      memory[11673] <=  254; /* free[253] */
      memory[11674] <=  255; /* free[254] */
      memory[11675] <=  256; /* free[255] */
      memory[11676] <=  257; /* free[256] */
      memory[11677] <=  258; /* free[257] */
      memory[11678] <=  259; /* free[258] */
      memory[11679] <=  260; /* free[259] */
      memory[11680] <=  261; /* free[260] */
      memory[11681] <=  262; /* free[261] */
      memory[11682] <=  263; /* free[262] */
      memory[11683] <=  264; /* free[263] */
      memory[11684] <=  265; /* free[264] */
      memory[11685] <=  266; /* free[265] */
      memory[11686] <=  267; /* free[266] */
      memory[11687] <=  268; /* free[267] */
      memory[11688] <=  269; /* free[268] */
      memory[11689] <=  270; /* free[269] */
      memory[11690] <=  271; /* free[270] */
      memory[11691] <=  272; /* free[271] */
      memory[11692] <=  273; /* free[272] */
      memory[11693] <=  274; /* free[273] */
      memory[11694] <=  275; /* free[274] */
      memory[11695] <=  276; /* free[275] */
      memory[11696] <=  277; /* free[276] */
      memory[11697] <=  278; /* free[277] */
      memory[11698] <=  279; /* free[278] */
      memory[11699] <=  280; /* free[279] */
      memory[11700] <=  281; /* free[280] */
      memory[11701] <=  282; /* free[281] */
      memory[11702] <=  283; /* free[282] */
      memory[11703] <=  284; /* free[283] */
      memory[11704] <=  285; /* free[284] */
      memory[11705] <=  286; /* free[285] */
      memory[11706] <=  287; /* free[286] */
      memory[11707] <=  288; /* free[287] */
      memory[11708] <=  289; /* free[288] */
      memory[11709] <=  290; /* free[289] */
      memory[11710] <=  291; /* free[290] */
      memory[11711] <=  292; /* free[291] */
      memory[11712] <=  293; /* free[292] */
      memory[11713] <=  294; /* free[293] */
      memory[11714] <=  295; /* free[294] */
      memory[11715] <=  296; /* free[295] */
      memory[11716] <=  297; /* free[296] */
      memory[11717] <=  298; /* free[297] */
      memory[11718] <=  299; /* free[298] */
      memory[11719] <=  300; /* free[299] */
      memory[11720] <=  301; /* free[300] */
      memory[11721] <=  302; /* free[301] */
      memory[11722] <=  303; /* free[302] */
      memory[11723] <=  304; /* free[303] */
      memory[11724] <=  305; /* free[304] */
      memory[11725] <=  306; /* free[305] */
      memory[11726] <=  307; /* free[306] */
      memory[11727] <=  308; /* free[307] */
      memory[11728] <=  309; /* free[308] */
      memory[11729] <=  310; /* free[309] */
      memory[11730] <=  311; /* free[310] */
      memory[11731] <=  312; /* free[311] */
      memory[11732] <=  313; /* free[312] */
      memory[11733] <=  314; /* free[313] */
      memory[11734] <=  315; /* free[314] */
      memory[11735] <=  316; /* free[315] */
      memory[11736] <=  317; /* free[316] */
      memory[11737] <=  318; /* free[317] */
      memory[11738] <=  319; /* free[318] */
      memory[11739] <=  320; /* free[319] */
      memory[11740] <=  321; /* free[320] */
      memory[11741] <=  322; /* free[321] */
      memory[11742] <=  323; /* free[322] */
      memory[11743] <=  324; /* free[323] */
      memory[11744] <=  325; /* free[324] */
      memory[11745] <=  326; /* free[325] */
      memory[11746] <=  327; /* free[326] */
      memory[11747] <=  328; /* free[327] */
      memory[11748] <=  329; /* free[328] */
      memory[11749] <=  330; /* free[329] */
      memory[11750] <=  331; /* free[330] */
      memory[11751] <=  332; /* free[331] */
      memory[11752] <=  333; /* free[332] */
      memory[11753] <=  334; /* free[333] */
      memory[11754] <=  335; /* free[334] */
      memory[11755] <=  336; /* free[335] */
      memory[11756] <=  337; /* free[336] */
      memory[11757] <=  338; /* free[337] */
      memory[11758] <=  339; /* free[338] */
      memory[11759] <=  340; /* free[339] */
      memory[11760] <=  341; /* free[340] */
      memory[11761] <=  342; /* free[341] */
      memory[11762] <=  343; /* free[342] */
      memory[11763] <=  344; /* free[343] */
      memory[11764] <=  345; /* free[344] */
      memory[11765] <=  346; /* free[345] */
      memory[11766] <=  347; /* free[346] */
      memory[11767] <=  348; /* free[347] */
      memory[11768] <=  349; /* free[348] */
      memory[11769] <=  350; /* free[349] */
      memory[11770] <=  351; /* free[350] */
      memory[11771] <=  352; /* free[351] */
      memory[11772] <=  353; /* free[352] */
      memory[11773] <=  354; /* free[353] */
      memory[11774] <=  355; /* free[354] */
      memory[11775] <=  356; /* free[355] */
      memory[11776] <=  357; /* free[356] */
      memory[11777] <=  358; /* free[357] */
      memory[11778] <=  359; /* free[358] */
      memory[11779] <=  360; /* free[359] */
      memory[11780] <=  361; /* free[360] */
      memory[11781] <=  362; /* free[361] */
      memory[11782] <=  363; /* free[362] */
      memory[11783] <=  364; /* free[363] */
      memory[11784] <=  365; /* free[364] */
      memory[11785] <=  366; /* free[365] */
      memory[11786] <=  367; /* free[366] */
      memory[11787] <=  368; /* free[367] */
      memory[11788] <=  369; /* free[368] */
      memory[11789] <=  370; /* free[369] */
      memory[11790] <=  371; /* free[370] */
      memory[11791] <=  372; /* free[371] */
      memory[11792] <=  373; /* free[372] */
      memory[11793] <=  374; /* free[373] */
      memory[11794] <=  375; /* free[374] */
      memory[11795] <=  376; /* free[375] */
      memory[11796] <=  377; /* free[376] */
      memory[11797] <=  378; /* free[377] */
      memory[11798] <=  379; /* free[378] */
      memory[11799] <=  380; /* free[379] */
      memory[11800] <=  381; /* free[380] */
      memory[11801] <=  382; /* free[381] */
      memory[11802] <=  383; /* free[382] */
      memory[11803] <=  384; /* free[383] */
      memory[11804] <=  385; /* free[384] */
      memory[11805] <=  386; /* free[385] */
      memory[11806] <=  387; /* free[386] */
      memory[11807] <=  388; /* free[387] */
      memory[11808] <=  389; /* free[388] */
      memory[11809] <=  390; /* free[389] */
      memory[11810] <=  391; /* free[390] */
      memory[11811] <=  392; /* free[391] */
      memory[11812] <=  393; /* free[392] */
      memory[11813] <=  394; /* free[393] */
      memory[11814] <=  395; /* free[394] */
      memory[11815] <=  396; /* free[395] */
      memory[11816] <=  397; /* free[396] */
      memory[11817] <=  398; /* free[397] */
      memory[11818] <=  399; /* free[398] */
      memory[11819] <=  400; /* free[399] */
      memory[11820] <=  401; /* free[400] */
      memory[11821] <=  402; /* free[401] */
      memory[11822] <=  403; /* free[402] */
      memory[11823] <=  404; /* free[403] */
      memory[11824] <=  405; /* free[404] */
      memory[11825] <=  406; /* free[405] */
      memory[11826] <=  407; /* free[406] */
      memory[11827] <=  408; /* free[407] */
      memory[11828] <=  409; /* free[408] */
      memory[11829] <=  410; /* free[409] */
      memory[11830] <=  411; /* free[410] */
      memory[11831] <=  412; /* free[411] */
      memory[11832] <=  413; /* free[412] */
      memory[11833] <=  414; /* free[413] */
      memory[11834] <=  415; /* free[414] */
      memory[11835] <=  416; /* free[415] */
      memory[11836] <=  417; /* free[416] */
      memory[11837] <=  418; /* free[417] */
      memory[11838] <=  419; /* free[418] */
      memory[11839] <=  420; /* free[419] */
      memory[11840] <=  421; /* free[420] */
      memory[11841] <=  422; /* free[421] */
      memory[11842] <=  423; /* free[422] */
      memory[11843] <=  424; /* free[423] */
      memory[11844] <=  425; /* free[424] */
      memory[11845] <=  426; /* free[425] */
      memory[11846] <=  427; /* free[426] */
      memory[11847] <=  428; /* free[427] */
      memory[11848] <=  429; /* free[428] */
      memory[11849] <=  430; /* free[429] */
      memory[11850] <=  431; /* free[430] */
      memory[11851] <=  432; /* free[431] */
      memory[11852] <=  433; /* free[432] */
      memory[11853] <=  434; /* free[433] */
      memory[11854] <=  435; /* free[434] */
      memory[11855] <=  436; /* free[435] */
      memory[11856] <=  437; /* free[436] */
      memory[11857] <=  438; /* free[437] */
      memory[11858] <=  439; /* free[438] */
      memory[11859] <=  440; /* free[439] */
      memory[11860] <=  441; /* free[440] */
      memory[11861] <=  442; /* free[441] */
      memory[11862] <=  443; /* free[442] */
      memory[11863] <=  444; /* free[443] */
      memory[11864] <=  445; /* free[444] */
      memory[11865] <=  446; /* free[445] */
      memory[11866] <=  447; /* free[446] */
      memory[11867] <=  448; /* free[447] */
      memory[11868] <=  449; /* free[448] */
      memory[11869] <=  450; /* free[449] */
      memory[11870] <=  451; /* free[450] */
      memory[11871] <=  452; /* free[451] */
      memory[11872] <=  453; /* free[452] */
      memory[11873] <=  454; /* free[453] */
      memory[11874] <=  455; /* free[454] */
      memory[11875] <=  456; /* free[455] */
      memory[11876] <=  457; /* free[456] */
      memory[11877] <=  458; /* free[457] */
      memory[11878] <=  459; /* free[458] */
      memory[11879] <=  460; /* free[459] */
      memory[11880] <=  461; /* free[460] */
      memory[11881] <=  462; /* free[461] */
      memory[11882] <=  463; /* free[462] */
      memory[11883] <=  464; /* free[463] */
      memory[11884] <=  465; /* free[464] */
      memory[11885] <=  466; /* free[465] */
      memory[11886] <=  467; /* free[466] */
      memory[11887] <=  468; /* free[467] */
      memory[11888] <=  469; /* free[468] */
      memory[11889] <=  470; /* free[469] */
      memory[11890] <=  471; /* free[470] */
      memory[11891] <=  472; /* free[471] */
      memory[11892] <=  473; /* free[472] */
      memory[11893] <=  474; /* free[473] */
      memory[11894] <=  475; /* free[474] */
      memory[11895] <=  476; /* free[475] */
      memory[11896] <=  477; /* free[476] */
      memory[11897] <=  478; /* free[477] */
      memory[11898] <=  479; /* free[478] */
      memory[11899] <=  480; /* free[479] */
      memory[11900] <=  481; /* free[480] */
      memory[11901] <=  482; /* free[481] */
      memory[11902] <=  483; /* free[482] */
      memory[11903] <=  484; /* free[483] */
      memory[11904] <=  485; /* free[484] */
      memory[11905] <=  486; /* free[485] */
      memory[11906] <=  487; /* free[486] */
      memory[11907] <=  488; /* free[487] */
      memory[11908] <=  489; /* free[488] */
      memory[11909] <=  490; /* free[489] */
      memory[11910] <=  491; /* free[490] */
      memory[11911] <=  492; /* free[491] */
      memory[11912] <=  493; /* free[492] */
      memory[11913] <=  494; /* free[493] */
      memory[11914] <=  495; /* free[494] */
      memory[11915] <=  496; /* free[495] */
      memory[11916] <=  497; /* free[496] */
      memory[11917] <=  498; /* free[497] */
      memory[11918] <=  499; /* free[498] */
      memory[11919] <=  500; /* free[499] */
      memory[11920] <=  501; /* free[500] */
      memory[11921] <=  502; /* free[501] */
      memory[11922] <=  503; /* free[502] */
      memory[11923] <=  504; /* free[503] */
      memory[11924] <=  505; /* free[504] */
      memory[11925] <=  506; /* free[505] */
      memory[11926] <=  507; /* free[506] */
      memory[11927] <=  508; /* free[507] */
      memory[11928] <=  509; /* free[508] */
      memory[11929] <=  510; /* free[509] */
      memory[11930] <=  511; /* free[510] */
      memory[11931] <=  512; /* free[511] */
      memory[11932] <=  513; /* free[512] */
      memory[11933] <=  514; /* free[513] */
      memory[11934] <=  515; /* free[514] */
      memory[11935] <=  516; /* free[515] */
      memory[11936] <=  517; /* free[516] */
      memory[11937] <=  518; /* free[517] */
      memory[11938] <=  519; /* free[518] */
      memory[11939] <=  520; /* free[519] */
      memory[11940] <=  521; /* free[520] */
      memory[11941] <=  522; /* free[521] */
      memory[11942] <=  523; /* free[522] */
      memory[11943] <=  524; /* free[523] */
      memory[11944] <=  525; /* free[524] */
      memory[11945] <=  526; /* free[525] */
      memory[11946] <=  527; /* free[526] */
      memory[11947] <=  528; /* free[527] */
      memory[11948] <=  529; /* free[528] */
      memory[11949] <=  530; /* free[529] */
      memory[11950] <=  531; /* free[530] */
      memory[11951] <=  532; /* free[531] */
      memory[11952] <=  533; /* free[532] */
      memory[11953] <=  534; /* free[533] */
      memory[11954] <=  535; /* free[534] */
      memory[11955] <=  536; /* free[535] */
      memory[11956] <=  537; /* free[536] */
      memory[11957] <=  538; /* free[537] */
      memory[11958] <=  539; /* free[538] */
      memory[11959] <=  540; /* free[539] */
      memory[11960] <=  541; /* free[540] */
      memory[11961] <=  542; /* free[541] */
      memory[11962] <=  543; /* free[542] */
      memory[11963] <=  544; /* free[543] */
      memory[11964] <=  545; /* free[544] */
      memory[11965] <=  546; /* free[545] */
      memory[11966] <=  547; /* free[546] */
      memory[11967] <=  548; /* free[547] */
      memory[11968] <=  549; /* free[548] */
      memory[11969] <=  550; /* free[549] */
      memory[11970] <=  551; /* free[550] */
      memory[11971] <=  552; /* free[551] */
      memory[11972] <=  553; /* free[552] */
      memory[11973] <=  554; /* free[553] */
      memory[11974] <=  555; /* free[554] */
      memory[11975] <=  556; /* free[555] */
      memory[11976] <=  557; /* free[556] */
      memory[11977] <=  558; /* free[557] */
      memory[11978] <=  559; /* free[558] */
      memory[11979] <=  560; /* free[559] */
      memory[11980] <=  561; /* free[560] */
      memory[11981] <=  562; /* free[561] */
      memory[11982] <=  563; /* free[562] */
      memory[11983] <=  564; /* free[563] */
      memory[11984] <=  565; /* free[564] */
      memory[11985] <=  566; /* free[565] */
      memory[11986] <=  567; /* free[566] */
      memory[11987] <=  568; /* free[567] */
      memory[11988] <=  569; /* free[568] */
      memory[11989] <=  570; /* free[569] */
      memory[11990] <=  571; /* free[570] */
      memory[11991] <=  572; /* free[571] */
      memory[11992] <=  573; /* free[572] */
      memory[11993] <=  574; /* free[573] */
      memory[11994] <=  575; /* free[574] */
      memory[11995] <=  576; /* free[575] */
      memory[11996] <=  577; /* free[576] */
      memory[11997] <=  578; /* free[577] */
      memory[11998] <=  579; /* free[578] */
      memory[11999] <=  580; /* free[579] */
      memory[12000] <=  581; /* free[580] */
      memory[12001] <=  582; /* free[581] */
      memory[12002] <=  583; /* free[582] */
      memory[12003] <=  584; /* free[583] */
      memory[12004] <=  585; /* free[584] */
      memory[12005] <=  586; /* free[585] */
      memory[12006] <=  587; /* free[586] */
      memory[12007] <=  588; /* free[587] */
      memory[12008] <=  589; /* free[588] */
      memory[12009] <=  590; /* free[589] */
      memory[12010] <=  591; /* free[590] */
      memory[12011] <=  592; /* free[591] */
      memory[12012] <=  593; /* free[592] */
      memory[12013] <=  594; /* free[593] */
      memory[12014] <=  595; /* free[594] */
      memory[12015] <=  596; /* free[595] */
      memory[12016] <=  597; /* free[596] */
      memory[12017] <=  598; /* free[597] */
      memory[12018] <=  599; /* free[598] */
      memory[12020] <=    1; /* f_success */
      memory[12021] <=    1; /* hasLeavesForChildren */
      memory[12022] <=    1; /* isALeaf */
      memory[12026] <=    1; /* isLeaf[1] */
      memory[12027] <=    1; /* isLeaf[2] */
      memory[12028] <=    1; /* isLeaf[3] */
      memory[12029] <=    1; /* isLeaf[4] */
      memory[12030] <=    1; /* isLeaf[5] */
      memory[12031] <=    1; /* isLeaf[6] */
      memory[12032] <=    1; /* isLeaf[7] */
      memory[12033] <=    1; /* isLeaf[8] */
      memory[12034] <=    1; /* isLeaf[9] */
      memory[12035] <=    1; /* isLeaf[10] */
      memory[12036] <=    1; /* isLeaf[11] */
      memory[12037] <=    1; /* isLeaf[12] */
      memory[12038] <=    1; /* isLeaf[13] */
      memory[12039] <=    1; /* isLeaf[14] */
      memory[12040] <=    1; /* isLeaf[15] */
      memory[12041] <=    1; /* isLeaf[16] */
      memory[12042] <=   -1; /* isLeaf[17] */
      memory[12626] <=   16; /* keys[0,0] */
      memory[12627] <=   32; /* keys[0,1] */
      memory[12628] <=   48; /* keys[0,2] */
      memory[12629] <=   64; /* keys[0,3] */
      memory[12630] <=   80; /* keys[0,4] */
      memory[12631] <=   96; /* keys[0,5] */
      memory[12632] <=  112; /* keys[0,6] */
      memory[12633] <=  128; /* keys[0,7] */
      memory[12634] <=  144; /* keys[0,8] */
      memory[12635] <=  160; /* keys[0,9] */
      memory[12636] <=  176; /* keys[0,10] */
      memory[12637] <=  192; /* keys[0,11] */
      memory[12638] <=  208; /* keys[0,12] */
      memory[12639] <=  224; /* keys[0,13] */
      memory[12640] <=  240; /* keys[0,14] */
      memory[12644] <=    1; /* keys[1,0] */
      memory[12645] <=    2; /* keys[1,1] */
      memory[12646] <=    3; /* keys[1,2] */
      memory[12647] <=    4; /* keys[1,3] */
      memory[12648] <=    5; /* keys[1,4] */
      memory[12649] <=    6; /* keys[1,5] */
      memory[12650] <=    7; /* keys[1,6] */
      memory[12651] <=    8; /* keys[1,7] */
      memory[12652] <=    9; /* keys[1,8] */
      memory[12653] <=   10; /* keys[1,9] */
      memory[12654] <=   11; /* keys[1,10] */
      memory[12655] <=   12; /* keys[1,11] */
      memory[12656] <=   13; /* keys[1,12] */
      memory[12657] <=   14; /* keys[1,13] */
      memory[12658] <=   15; /* keys[1,14] */
      memory[12659] <=   16; /* keys[1,15] */
      memory[12662] <=  241; /* keys[2,0] */
      memory[12663] <=  242; /* keys[2,1] */
      memory[12664] <=  243; /* keys[2,2] */
      memory[12665] <=  244; /* keys[2,3] */
      memory[12666] <=  245; /* keys[2,4] */
      memory[12667] <=  246; /* keys[2,5] */
      memory[12668] <=  247; /* keys[2,6] */
      memory[12669] <=  248; /* keys[2,7] */
      memory[12670] <=  249; /* keys[2,8] */
      memory[12671] <=  250; /* keys[2,9] */
      memory[12672] <=  251; /* keys[2,10] */
      memory[12673] <=  252; /* keys[2,11] */
      memory[12674] <=  253; /* keys[2,12] */
      memory[12675] <=  254; /* keys[2,13] */
      memory[12676] <=  255; /* keys[2,14] */
      memory[12677] <=  256; /* keys[2,15] */
      memory[12680] <=   17; /* keys[3,0] */
      memory[12681] <=   18; /* keys[3,1] */
      memory[12682] <=   19; /* keys[3,2] */
      memory[12683] <=   20; /* keys[3,3] */
      memory[12684] <=   21; /* keys[3,4] */
      memory[12685] <=   22; /* keys[3,5] */
      memory[12686] <=   23; /* keys[3,6] */
      memory[12687] <=   24; /* keys[3,7] */
      memory[12688] <=   25; /* keys[3,8] */
      memory[12689] <=   26; /* keys[3,9] */
      memory[12690] <=   27; /* keys[3,10] */
      memory[12691] <=   28; /* keys[3,11] */
      memory[12692] <=   29; /* keys[3,12] */
      memory[12693] <=   30; /* keys[3,13] */
      memory[12694] <=   31; /* keys[3,14] */
      memory[12695] <=   32; /* keys[3,15] */
      memory[12698] <=   33; /* keys[4,0] */
      memory[12699] <=   34; /* keys[4,1] */
      memory[12700] <=   35; /* keys[4,2] */
      memory[12701] <=   36; /* keys[4,3] */
      memory[12702] <=   37; /* keys[4,4] */
      memory[12703] <=   38; /* keys[4,5] */
      memory[12704] <=   39; /* keys[4,6] */
      memory[12705] <=   40; /* keys[4,7] */
      memory[12706] <=   41; /* keys[4,8] */
      memory[12707] <=   42; /* keys[4,9] */
      memory[12708] <=   43; /* keys[4,10] */
      memory[12709] <=   44; /* keys[4,11] */
      memory[12710] <=   45; /* keys[4,12] */
      memory[12711] <=   46; /* keys[4,13] */
      memory[12712] <=   47; /* keys[4,14] */
      memory[12713] <=   48; /* keys[4,15] */
      memory[12716] <=   49; /* keys[5,0] */
      memory[12717] <=   50; /* keys[5,1] */
      memory[12718] <=   51; /* keys[5,2] */
      memory[12719] <=   52; /* keys[5,3] */
      memory[12720] <=   53; /* keys[5,4] */
      memory[12721] <=   54; /* keys[5,5] */
      memory[12722] <=   55; /* keys[5,6] */
      memory[12723] <=   56; /* keys[5,7] */
      memory[12724] <=   57; /* keys[5,8] */
      memory[12725] <=   58; /* keys[5,9] */
      memory[12726] <=   59; /* keys[5,10] */
      memory[12727] <=   60; /* keys[5,11] */
      memory[12728] <=   61; /* keys[5,12] */
      memory[12729] <=   62; /* keys[5,13] */
      memory[12730] <=   63; /* keys[5,14] */
      memory[12731] <=   64; /* keys[5,15] */
      memory[12734] <=   65; /* keys[6,0] */
      memory[12735] <=   66; /* keys[6,1] */
      memory[12736] <=   67; /* keys[6,2] */
      memory[12737] <=   68; /* keys[6,3] */
      memory[12738] <=   69; /* keys[6,4] */
      memory[12739] <=   70; /* keys[6,5] */
      memory[12740] <=   71; /* keys[6,6] */
      memory[12741] <=   72; /* keys[6,7] */
      memory[12742] <=   73; /* keys[6,8] */
      memory[12743] <=   74; /* keys[6,9] */
      memory[12744] <=   75; /* keys[6,10] */
      memory[12745] <=   76; /* keys[6,11] */
      memory[12746] <=   77; /* keys[6,12] */
      memory[12747] <=   78; /* keys[6,13] */
      memory[12748] <=   79; /* keys[6,14] */
      memory[12749] <=   80; /* keys[6,15] */
      memory[12752] <=   81; /* keys[7,0] */
      memory[12753] <=   82; /* keys[7,1] */
      memory[12754] <=   83; /* keys[7,2] */
      memory[12755] <=   84; /* keys[7,3] */
      memory[12756] <=   85; /* keys[7,4] */
      memory[12757] <=   86; /* keys[7,5] */
      memory[12758] <=   87; /* keys[7,6] */
      memory[12759] <=   88; /* keys[7,7] */
      memory[12760] <=   89; /* keys[7,8] */
      memory[12761] <=   90; /* keys[7,9] */
      memory[12762] <=   91; /* keys[7,10] */
      memory[12763] <=   92; /* keys[7,11] */
      memory[12764] <=   93; /* keys[7,12] */
      memory[12765] <=   94; /* keys[7,13] */
      memory[12766] <=   95; /* keys[7,14] */
      memory[12767] <=   96; /* keys[7,15] */
      memory[12770] <=   97; /* keys[8,0] */
      memory[12771] <=   98; /* keys[8,1] */
      memory[12772] <=   99; /* keys[8,2] */
      memory[12773] <=  100; /* keys[8,3] */
      memory[12774] <=  101; /* keys[8,4] */
      memory[12775] <=  102; /* keys[8,5] */
      memory[12776] <=  103; /* keys[8,6] */
      memory[12777] <=  104; /* keys[8,7] */
      memory[12778] <=  105; /* keys[8,8] */
      memory[12779] <=  106; /* keys[8,9] */
      memory[12780] <=  107; /* keys[8,10] */
      memory[12781] <=  108; /* keys[8,11] */
      memory[12782] <=  109; /* keys[8,12] */
      memory[12783] <=  110; /* keys[8,13] */
      memory[12784] <=  111; /* keys[8,14] */
      memory[12785] <=  112; /* keys[8,15] */
      memory[12788] <=  113; /* keys[9,0] */
      memory[12789] <=  114; /* keys[9,1] */
      memory[12790] <=  115; /* keys[9,2] */
      memory[12791] <=  116; /* keys[9,3] */
      memory[12792] <=  117; /* keys[9,4] */
      memory[12793] <=  118; /* keys[9,5] */
      memory[12794] <=  119; /* keys[9,6] */
      memory[12795] <=  120; /* keys[9,7] */
      memory[12796] <=  121; /* keys[9,8] */
      memory[12797] <=  122; /* keys[9,9] */
      memory[12798] <=  123; /* keys[9,10] */
      memory[12799] <=  124; /* keys[9,11] */
      memory[12800] <=  125; /* keys[9,12] */
      memory[12801] <=  126; /* keys[9,13] */
      memory[12802] <=  127; /* keys[9,14] */
      memory[12803] <=  128; /* keys[9,15] */
      memory[12806] <=  129; /* keys[10,0] */
      memory[12807] <=  130; /* keys[10,1] */
      memory[12808] <=  131; /* keys[10,2] */
      memory[12809] <=  132; /* keys[10,3] */
      memory[12810] <=  133; /* keys[10,4] */
      memory[12811] <=  134; /* keys[10,5] */
      memory[12812] <=  135; /* keys[10,6] */
      memory[12813] <=  136; /* keys[10,7] */
      memory[12814] <=  137; /* keys[10,8] */
      memory[12815] <=  138; /* keys[10,9] */
      memory[12816] <=  139; /* keys[10,10] */
      memory[12817] <=  140; /* keys[10,11] */
      memory[12818] <=  141; /* keys[10,12] */
      memory[12819] <=  142; /* keys[10,13] */
      memory[12820] <=  143; /* keys[10,14] */
      memory[12821] <=  144; /* keys[10,15] */
      memory[12824] <=  145; /* keys[11,0] */
      memory[12825] <=  146; /* keys[11,1] */
      memory[12826] <=  147; /* keys[11,2] */
      memory[12827] <=  148; /* keys[11,3] */
      memory[12828] <=  149; /* keys[11,4] */
      memory[12829] <=  150; /* keys[11,5] */
      memory[12830] <=  151; /* keys[11,6] */
      memory[12831] <=  152; /* keys[11,7] */
      memory[12832] <=  153; /* keys[11,8] */
      memory[12833] <=  154; /* keys[11,9] */
      memory[12834] <=  155; /* keys[11,10] */
      memory[12835] <=  156; /* keys[11,11] */
      memory[12836] <=  157; /* keys[11,12] */
      memory[12837] <=  158; /* keys[11,13] */
      memory[12838] <=  159; /* keys[11,14] */
      memory[12839] <=  160; /* keys[11,15] */
      memory[12842] <=  161; /* keys[12,0] */
      memory[12843] <=  162; /* keys[12,1] */
      memory[12844] <=  163; /* keys[12,2] */
      memory[12845] <=  164; /* keys[12,3] */
      memory[12846] <=  165; /* keys[12,4] */
      memory[12847] <=  166; /* keys[12,5] */
      memory[12848] <=  167; /* keys[12,6] */
      memory[12849] <=  168; /* keys[12,7] */
      memory[12850] <=  169; /* keys[12,8] */
      memory[12851] <=  170; /* keys[12,9] */
      memory[12852] <=  171; /* keys[12,10] */
      memory[12853] <=  172; /* keys[12,11] */
      memory[12854] <=  173; /* keys[12,12] */
      memory[12855] <=  174; /* keys[12,13] */
      memory[12856] <=  175; /* keys[12,14] */
      memory[12857] <=  176; /* keys[12,15] */
      memory[12860] <=  177; /* keys[13,0] */
      memory[12861] <=  178; /* keys[13,1] */
      memory[12862] <=  179; /* keys[13,2] */
      memory[12863] <=  180; /* keys[13,3] */
      memory[12864] <=  181; /* keys[13,4] */
      memory[12865] <=  182; /* keys[13,5] */
      memory[12866] <=  183; /* keys[13,6] */
      memory[12867] <=  184; /* keys[13,7] */
      memory[12868] <=  185; /* keys[13,8] */
      memory[12869] <=  186; /* keys[13,9] */
      memory[12870] <=  187; /* keys[13,10] */
      memory[12871] <=  188; /* keys[13,11] */
      memory[12872] <=  189; /* keys[13,12] */
      memory[12873] <=  190; /* keys[13,13] */
      memory[12874] <=  191; /* keys[13,14] */
      memory[12875] <=  192; /* keys[13,15] */
      memory[12878] <=  193; /* keys[14,0] */
      memory[12879] <=  194; /* keys[14,1] */
      memory[12880] <=  195; /* keys[14,2] */
      memory[12881] <=  196; /* keys[14,3] */
      memory[12882] <=  197; /* keys[14,4] */
      memory[12883] <=  198; /* keys[14,5] */
      memory[12884] <=  199; /* keys[14,6] */
      memory[12885] <=  200; /* keys[14,7] */
      memory[12886] <=  201; /* keys[14,8] */
      memory[12887] <=  202; /* keys[14,9] */
      memory[12888] <=  203; /* keys[14,10] */
      memory[12889] <=  204; /* keys[14,11] */
      memory[12890] <=  205; /* keys[14,12] */
      memory[12891] <=  206; /* keys[14,13] */
      memory[12892] <=  207; /* keys[14,14] */
      memory[12893] <=  208; /* keys[14,15] */
      memory[12896] <=  209; /* keys[15,0] */
      memory[12897] <=  210; /* keys[15,1] */
      memory[12898] <=  211; /* keys[15,2] */
      memory[12899] <=  212; /* keys[15,3] */
      memory[12900] <=  213; /* keys[15,4] */
      memory[12901] <=  214; /* keys[15,5] */
      memory[12902] <=  215; /* keys[15,6] */
      memory[12903] <=  216; /* keys[15,7] */
      memory[12904] <=  217; /* keys[15,8] */
      memory[12905] <=  218; /* keys[15,9] */
      memory[12906] <=  219; /* keys[15,10] */
      memory[12907] <=  220; /* keys[15,11] */
      memory[12908] <=  221; /* keys[15,12] */
      memory[12909] <=  222; /* keys[15,13] */
      memory[12910] <=  223; /* keys[15,14] */
      memory[12911] <=  224; /* keys[15,15] */
      memory[12914] <=  225; /* keys[16,0] */
      memory[12915] <=  226; /* keys[16,1] */
      memory[12916] <=  227; /* keys[16,2] */
      memory[12917] <=  228; /* keys[16,3] */
      memory[12918] <=  229; /* keys[16,4] */
      memory[12919] <=  230; /* keys[16,5] */
      memory[12920] <=  231; /* keys[16,6] */
      memory[12921] <=  232; /* keys[16,7] */
      memory[12922] <=  233; /* keys[16,8] */
      memory[12923] <=  234; /* keys[16,9] */
      memory[12924] <=  235; /* keys[16,10] */
      memory[12925] <=  236; /* keys[16,11] */
      memory[12926] <=  237; /* keys[16,12] */
      memory[12927] <=  238; /* keys[16,13] */
      memory[12928] <=  239; /* keys[16,14] */
      memory[12929] <=  240; /* keys[16,15] */
      memory[12932] <=   -1; /* keys[17,0] */
      memory[12933] <=   -1; /* keys[17,1] */
      memory[12934] <=   -1; /* keys[17,2] */
      memory[12935] <=   -1; /* keys[17,3] */
      memory[12936] <=   -1; /* keys[17,4] */
      memory[12937] <=   -1; /* keys[17,5] */
      memory[12938] <=   -1; /* keys[17,6] */
      memory[12939] <=   -1; /* keys[17,7] */
      memory[12940] <=   -1; /* keys[17,8] */
      memory[12941] <=   -1; /* keys[17,9] */
      memory[12942] <=   -1; /* keys[17,10] */
      memory[12943] <=   -1; /* keys[17,11] */
      memory[12944] <=   -1; /* keys[17,12] */
      memory[12945] <=   -1; /* keys[17,13] */
      memory[12946] <=   -1; /* keys[17,14] */
      memory[12947] <=   -1; /* keys[17,15] */
      memory[12948] <=   -1; /* keys[17,16] */
      memory[12949] <=   -1; /* keys[17,17] */
      memory[23426] <=   15; /* leafSize */
      memory[23427] <=   17; /* merge_indexLimit */
      memory[23428] <=   17; /* merge_indices */
      memory[23429] <=  249; /* merge_Key */
      memory[23430] <=   15; /* mergeLeftSibling_bs */
      memory[23431] <=   16; /* mergeLeftSibling_index */
      memory[23432] <=   15; /* mergeLeftSibling_l */
      memory[23433] <=   16; /* mergeLeftSibling_nl */
      memory[23434] <=   24; /* mergeLeftSibling_nlr */
      memory[23435] <=    8; /* mergeLeftSibling_nr */
      memory[23437] <=   16; /* mergeLeftSibling_r */
      memory[23441] <=    1; /* merge_loop */
      memory[23442] <=   15; /* mergeRightSibling_bs */
      memory[23444] <=   16; /* mergeRightSibling_index */
      memory[23446] <=   16; /* mergeRightSibling_l */
      memory[23447] <=    8; /* mergeRightSibling_nl */
      memory[23448] <=   16; /* mergeRightSibling_nlr */
      memory[23449] <=    8; /* mergeRightSibling_nr */
      memory[23451] <=  240; /* mergeRightSibling_pk */
      memory[23452] <=   17; /* mergeRightSibling_r */
      memory[23453] <=    8; /* mergeRightSibling_size */
      memory[23459] <=   16; /* mergeRoot_nP */
      memory[23464] <=    1; /* put_Data */
      memory[23465] <=  256; /* put_Key */
      memory[23469] <=    1; /* s_data */
      memory[23471] <=   17; /* setLeaf */
      memory[23473] <=   15; /* s_index */
      memory[23474] <=  256; /* s_key */
      memory[23483] <=  241; /* splitLeaf_F */
      memory[23484] <=  240; /* splitLeaf_fl */
      memory[23485] <=   15; /* splitLeaf_index */
      memory[23486] <=  240; /* splitLeaf_L */
      memory[23487] <=   17; /* splitLeaf_l */
      memory[23488] <=    2; /* splitLeaf_node */
      memory[23490] <=    9; /* splitLeafRoot_first */
      memory[23492] <=    8; /* splitLeafRoot_kv */
      memory[23493] <=    8; /* splitLeafRoot_last */
      memory[23494] <=    1; /* splitLeafRoot_l */
      memory[23495] <=    2; /* splitLeafRoot_r */
      memory[23518] <=   14; /* stuckInsertElementAt_I */
      memory[23519] <=   15; /* stuckInsertElementAt_i */
      memory[23520] <=   15; /* stuckInsertElementAt_L */
      memory[23521] <=   17; /* stuckRemoveElementAt_I */
      memory[23522] <=   16; /* stuckRemoveElementAt_i */
      memory[23523] <=   17; /* stuckRemoveElementAt_N */
      memory[23524] <=   15; /* stuckSearch_N */
      memory[23526] <=    1; /* stuckShift_I */
      memory[23527] <=    1; /* stuckShift_N */
      memory[23528] <=    2; /* stuck */

      memory[11413] <= 22; /* find key */

    end
    else begin                                                                  // Run
      //$display("%4d %4d %4d s=%4d f=%4d d=%4d", steps, step, intermediateValue, stop, found, data);
      case(step)
         0: begin intermediateValue <= memory[12025+memory[23467]/*root*/]/*isLeaf[root]*/; /* get 2 */ step <= step + 1; end
         1: begin memory[23468]/*rootIsLeaf*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         2: begin intermediateValue <= memory[23468]/*rootIsLeaf*/; /* get 1 */ step <= step + 1; end
         3: begin if (intermediateValue == 0) step <=   38; else step = step + 1;/* endIfEq*/    end
         4: begin memory[23528]/*stuck*/ <= 0; /* set 1 */ step <= step + 1; end
         5: begin intermediateValue <= memory[11413]/*find_Key*/; /* get 1 */ step <= step + 1; end
         6: begin memory[23474]/*s_key*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
         7: begin memory[23472]/*s_found*/ <= 0; /* set 1 */ step <= step + 1; end
         8: begin memory[23473]/*s_index*/ <= 0; /* set 1 */ step <= step + 1; end
         9: begin intermediateValue <= memory[5+memory[23528]/*stuck*/]/*current_size[stuck]*/; /* get 2 */ step <= step + 1; end
        10: begin memory[23524]/*stuckSearch_N*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        11: begin intermediateValue <= memory[23473]/*s_index*/ < memory[23524]/*stuckSearch_N*/ ? -1 : memory[23473]/*s_index*/ == memory[23524]/*stuckSearch_N*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
        12: begin if (intermediateValue >= 0) step <=   27; else step = step + 1;/* endIfGe*/    end
        13: begin intermediateValue <= memory[23474]/*s_key*/ < memory[12626+memory[23528]/*stuck*/*18+memory[23473]/*s_index*/]/*keys[s_index,stuck]*/ ? -1 : memory[23474]/*s_key*/ == memory[12626+memory[23528]/*stuck*/*18+memory[23473]/*s_index*/]/*keys[s_index,stuck]*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
        14: begin if (intermediateValue != 0) step <=   21; else step = step + 1;/* endIfNe*/    end
        15: begin memory[23472]/*s_found*/ <= 1; /* set 1 */ step <= step + 1; end
        16: begin intermediateValue <= memory[12626+memory[23528]/*stuck*/*18+memory[23473]/*s_index*/]/*keys[s_index,stuck]*/; /* get 3 */ step <= step + 1; end
        17: begin memory[23474]/*s_key*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        18: begin intermediateValue <= memory[605+memory[23528]/*stuck*/*18+memory[23473]/*s_index*/]/*data[s_index,stuck]*/; /* get 3 */ step <= step + 1; end
        19: begin memory[23469]/*s_data*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        20: begin step <=   27; /* end */ end
        21: begin intermediateValue <= memory[23473]/*s_index*/; /* get 1 */ step <= step + 1; end
        22: begin intermediateValue <= 1 + intermediateValue;  /* add 1 */ step <= step + 1; end
        23: begin memory[23473]/*s_index*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        24: begin intermediateValue <= memory[23473]/*s_index*/ < memory[23524]/*stuckSearch_N*/ ? -1 : memory[23473]/*s_index*/ == memory[23524]/*stuckSearch_N*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
        25: begin if (intermediateValue >= 0) step <=   27; else step = step + 1;/* endIfGe*/    end
        26: begin step <= 11; /* start */ end
        27: begin intermediateValue <= memory[23467]/*root*/; /* get 1 */ step <= step + 1; end
        28: begin memory[11418]/*f_leaf*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        29: begin intermediateValue <= memory[23472]/*s_found*/; /* get 1 */ step <= step + 1; end
        30: begin memory[11408]/*f_found*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        31: begin intermediateValue <= memory[23473]/*s_index*/; /* get 1 */ step <= step + 1; end
        32: begin memory[11412]/*f_index*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        33: begin intermediateValue <= memory[23474]/*s_key*/; /* get 1 */ step <= step + 1; end
        34: begin memory[11417]/*f_key*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        35: begin intermediateValue <= memory[23469]/*s_data*/; /* get 1 */ step <= step + 1; end
        36: begin memory[11407]/*f_data*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        37: begin step <=   127; /* end */ end
        38: begin intermediateValue <= memory[23467]/*root*/; /* get 1 */ step <= step + 1; end
        39: begin memory[23463]/*parent*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        40: begin memory[11414] <= 0; /* clear 1 */ step <= step + 1; end
        41: begin intermediateValue <= memory[23463]/*parent*/; /* get 1 */ step <= step + 1; end
        42: begin memory[23528]/*stuck*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        43: begin intermediateValue <= memory[11413]/*find_Key*/; /* get 1 */ step <= step + 1; end
        44: begin memory[23474]/*s_key*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        45: begin memory[23472]/*s_found*/ <= 0; /* set 1 */ step <= step + 1; end
        46: begin memory[23473]/*s_index*/ <= 0; /* set 1 */ step <= step + 1; end
        47: begin intermediateValue <= memory[5+memory[23528]/*stuck*/]/*current_size[stuck]*/; /* get 2 */ step <= step + 1; end
        48: begin memory[23524]/*stuckSearch_N*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        49: begin intermediateValue <= memory[23524]/*stuckSearch_N*/; /* get 1 */ step <= step + 1; end
        50: begin intermediateValue <= -1 + intermediateValue;  /* add 1 */ step <= step + 1; end
        51: begin memory[23524]/*stuckSearch_N*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        52: begin intermediateValue <= memory[23473]/*s_index*/ < memory[23524]/*stuckSearch_N*/ ? -1 : memory[23473]/*s_index*/ == memory[23524]/*stuckSearch_N*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
        53: begin if (intermediateValue >= 0) step <=   68; else step = step + 1;/* endIfGe*/    end
        54: begin intermediateValue <= memory[23474]/*s_key*/ < memory[12626+memory[23528]/*stuck*/*18+memory[23473]/*s_index*/]/*keys[s_index,stuck]*/ ? -1 : memory[23474]/*s_key*/ == memory[12626+memory[23528]/*stuck*/*18+memory[23473]/*s_index*/]/*keys[s_index,stuck]*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
        55: begin if (intermediateValue >  0) step <=   62; else step = step + 1;/* endIfGt*/    end
        56: begin memory[23472]/*s_found*/ <= 1; /* set 1 */ step <= step + 1; end
        57: begin intermediateValue <= memory[12626+memory[23528]/*stuck*/*18+memory[23473]/*s_index*/]/*keys[s_index,stuck]*/; /* get 3 */ step <= step + 1; end
        58: begin memory[23474]/*s_key*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        59: begin intermediateValue <= memory[605+memory[23528]/*stuck*/*18+memory[23473]/*s_index*/]/*data[s_index,stuck]*/; /* get 3 */ step <= step + 1; end
        60: begin memory[23469]/*s_data*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        61: begin step <=   68; /* end */ end
        62: begin intermediateValue <= memory[23473]/*s_index*/; /* get 1 */ step <= step + 1; end
        63: begin intermediateValue <= 1 + intermediateValue;  /* add 1 */ step <= step + 1; end
        64: begin memory[23473]/*s_index*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        65: begin intermediateValue <= memory[23473]/*s_index*/ < memory[23524]/*stuckSearch_N*/ ? -1 : memory[23473]/*s_index*/ == memory[23524]/*stuckSearch_N*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
        66: begin if (intermediateValue >= 0) step <=   68; else step = step + 1;/* endIfGe*/    end
        67: begin step <= 52; /* start */ end
        68: begin intermediateValue <= memory[12626+memory[23528]/*stuck*/*18+memory[23473]/*s_index*/]/*keys[s_index,stuck]*/; /* get 3 */ step <= step + 1; end
        69: begin memory[23474]/*s_key*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        70: begin intermediateValue <= memory[605+memory[23528]/*stuck*/*18+memory[23473]/*s_index*/]/*data[s_index,stuck]*/; /* get 3 */ step <= step + 1; end
        71: begin memory[23469]/*s_data*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        72: begin intermediateValue <= memory[23469]/*s_data*/; /* get 1 */ step <= step + 1; end
        73: begin memory[4]/*child*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        74: begin intermediateValue <= memory[4]/*child*/; /* get 1 */ step <= step + 1; end
        75: begin memory[12022]/*isALeaf*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        76: begin intermediateValue <= memory[12025+memory[12022]/*isALeaf*/]/*isLeaf[isALeaf]*/; /* get 2 */ step <= step + 1; end
        77: begin memory[12022]/*isALeaf*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        78: begin intermediateValue <= memory[12022]/*isALeaf*/; /* get 1 */ step <= step + 1; end
        79: begin if (intermediateValue == 0) step <=   117; else step = step + 1;/* endIfEq*/    end
        80: begin intermediateValue <= memory[4]/*child*/; /* get 1 */ step <= step + 1; end
        81: begin memory[23528]/*stuck*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        82: begin intermediateValue <= memory[11413]/*find_Key*/; /* get 1 */ step <= step + 1; end
        83: begin memory[23474]/*s_key*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        84: begin memory[23472]/*s_found*/ <= 0; /* set 1 */ step <= step + 1; end
        85: begin memory[23473]/*s_index*/ <= 0; /* set 1 */ step <= step + 1; end
        86: begin intermediateValue <= memory[5+memory[23528]/*stuck*/]/*current_size[stuck]*/; /* get 2 */ step <= step + 1; end
        87: begin memory[23524]/*stuckSearch_N*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        88: begin intermediateValue <= memory[23473]/*s_index*/ < memory[23524]/*stuckSearch_N*/ ? -1 : memory[23473]/*s_index*/ == memory[23524]/*stuckSearch_N*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
        89: begin if (intermediateValue >= 0) step <=   104; else step = step + 1;/* endIfGe*/    end
        90: begin intermediateValue <= memory[23474]/*s_key*/ < memory[12626+memory[23528]/*stuck*/*18+memory[23473]/*s_index*/]/*keys[s_index,stuck]*/ ? -1 : memory[23474]/*s_key*/ == memory[12626+memory[23528]/*stuck*/*18+memory[23473]/*s_index*/]/*keys[s_index,stuck]*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
        91: begin if (intermediateValue != 0) step <=   98; else step = step + 1;/* endIfNe*/    end
        92: begin memory[23472]/*s_found*/ <= 1; /* set 1 */ step <= step + 1; end
        93: begin intermediateValue <= memory[12626+memory[23528]/*stuck*/*18+memory[23473]/*s_index*/]/*keys[s_index,stuck]*/; /* get 3 */ step <= step + 1; end
        94: begin memory[23474]/*s_key*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        95: begin intermediateValue <= memory[605+memory[23528]/*stuck*/*18+memory[23473]/*s_index*/]/*data[s_index,stuck]*/; /* get 3 */ step <= step + 1; end
        96: begin memory[23469]/*s_data*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
        97: begin step <=   104; /* end */ end
        98: begin intermediateValue <= memory[23473]/*s_index*/; /* get 1 */ step <= step + 1; end
        99: begin intermediateValue <= 1 + intermediateValue;  /* add 1 */ step <= step + 1; end
       100: begin memory[23473]/*s_index*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
       101: begin intermediateValue <= memory[23473]/*s_index*/ < memory[23524]/*stuckSearch_N*/ ? -1 : memory[23473]/*s_index*/ == memory[23524]/*stuckSearch_N*/ ?  0 : +1; /* compare 2 */ step <= step + 1; end
       102: begin if (intermediateValue >= 0) step <=   104; else step = step + 1;/* endIfGe*/    end
       103: begin step <= 88; /* start */ end
       104: begin intermediateValue <= memory[4]/*child*/; /* get 1 */ step <= step + 1; end
       105: begin memory[11415]/*find_result_leaf*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
       106: begin intermediateValue <= memory[11415]/*find_result_leaf*/; /* get 1 */ step <= step + 1; end
       107: begin memory[11418]/*f_leaf*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
       108: begin intermediateValue <= memory[23472]/*s_found*/; /* get 1 */ step <= step + 1; end
       109: begin memory[11408]/*f_found*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
       110: begin intermediateValue <= memory[23473]/*s_index*/; /* get 1 */ step <= step + 1; end
       111: begin memory[11412]/*f_index*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
       112: begin intermediateValue <= memory[23474]/*s_key*/; /* get 1 */ step <= step + 1; end
       113: begin memory[11417]/*f_key*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
       114: begin intermediateValue <= memory[23469]/*s_data*/; /* get 1 */ step <= step + 1; end
       115: begin memory[11407]/*f_data*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
       116: begin step <=   127; /* end */ end
       117: begin intermediateValue <= memory[4]/*child*/; /* get 1 */ step <= step + 1; end
       118: begin memory[23463]/*parent*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
       119: begin intermediateValue <= memory[11414]/*find_loop*/; /* get 1 */ step <= step + 1; end
       120: begin intermediateValue <= 1 + intermediateValue;  /* add 1 */ step <= step + 1; end
       121: begin memory[11414]/*find_loop*/ <= intermediateValue; /* set 1 */ step <= step + 1; end
       122: begin intermediateValue <= memory[11414]/*find_loop*/; /* get 1 */ step <= step + 1; end
       123: begin intermediateValue <= 9 <  intermediateValue ? -1 : 9 == intermediateValue ?  0 : +1; /* compare 1 */ step <= step + 1; end
       124: begin if (intermediateValue >= 0) step <=   126; else step = step + 1;/* endIfGe*/    end
       125: begin step <= 41; /* start */ end
       126: begin stopped <= 1; end

        default: stopped <= 1;
      endcase
      steps    <= steps + 1;
    end // Execute
  end // Always
endmodule
